// This file contains sigmoid and sigmoid prime table
// These are NOT parameterized for bit widths because that's too complicated
// Original settings are given below. If other bit width settings are desired, change manually

/*  SIGMOID TABLE:
	Original z = 16b = 1,5,10 => -32 to +32
	Domain z used here = 10b = 1,3,6 => -8 to +8, 0.015625 precision. These are bits [13:4] of original z
	When z<-8, f(z)=0. When z>8, f(z)=1. When z=0, f(z)=0.5
	Range f(z) = 8b = 0,0,8 => 0 to 1, 0.00390625 precision.
	Final sigmoid output value = 16b = 1,5,10. 6 MSB and 2 LSB are all 0. Bits [9:2] of final value are calculated f(z) */
module sigmoid_t #(
	parameter width = 16, 
	parameter int_bits = 10,
	parameter frac_bits = 21
)(
	input clk,
	input [width-1:0] z, //1+5+10
	output reg [width-1:0] sigmoid_out //1+5+10
);
	
	reg [20:0] sigmoid; //calculated f(z)
/*
	real real_z, real_sigmoid;

	

	always @(posedge clk)begin
		real_z = z/2**(frac_bits)-z[width-1]*2.0**(1+int_bits);
		real_sigmoid = 1.0/(1+2.71828**(-real_z));
		sigmoid_out = real_sigmoid*2**(frac_bits);
	end*/

	always @(posedge clk)
		sigmoid_out = (z[width-1:width-int_bits+2] == 0 || (&z[width-1:width-int_bits+2] ))?
			{{(int_bits+1){1'b0}}, sigmoid}: 
			(z[width-1])?  1: {1'b1, {(frac_bits){1'b0}}}-1;
	// If condition is not met, z is too high or too low. In that case, f'(z)=0

	always @(z[frac_bits+4:frac_bits-9])
	case (z[frac_bits+4:frac_bits-9])

		//sign, 4bits_i, 10bits_f ~ 0.015625  --->   8bits_f ~ 0.00390625
		14'b10000000000000:	sigmoid = 21'b000000000000000000001;
		14'b10000000000001:	sigmoid = 21'b000000000000000000001;
		14'b10000000000010:	sigmoid = 21'b000000000000000000001;
		14'b10000000000011:	sigmoid = 21'b000000000000000000001;
		14'b10000000000100:	sigmoid = 21'b000000000000000000001;
		14'b10000000000101:	sigmoid = 21'b000000000000000000001;
		14'b10000000000110:	sigmoid = 21'b000000000000000000001;
		14'b10000000000111:	sigmoid = 21'b000000000000000000001;
		14'b10000000001000:	sigmoid = 21'b000000000000000000001;
		14'b10000000001001:	sigmoid = 21'b000000000000000000001;
		14'b10000000001010:	sigmoid = 21'b000000000000000000001;
		14'b10000000001011:	sigmoid = 21'b000000000000000000001;
		14'b10000000001100:	sigmoid = 21'b000000000000000000001;
		14'b10000000001101:	sigmoid = 21'b000000000000000000001;
		14'b10000000001110:	sigmoid = 21'b000000000000000000001;
		14'b10000000001111:	sigmoid = 21'b000000000000000000001;
		14'b10000000010000:	sigmoid = 21'b000000000000000000001;
		14'b10000000010001:	sigmoid = 21'b000000000000000000001;
		14'b10000000010010:	sigmoid = 21'b000000000000000000001;
		14'b10000000010011:	sigmoid = 21'b000000000000000000001;
		14'b10000000010100:	sigmoid = 21'b000000000000000000001;
		14'b10000000010101:	sigmoid = 21'b000000000000000000001;
		14'b10000000010110:	sigmoid = 21'b000000000000000000001;
		14'b10000000010111:	sigmoid = 21'b000000000000000000001;
		14'b10000000011000:	sigmoid = 21'b000000000000000000001;
		14'b10000000011001:	sigmoid = 21'b000000000000000000001;
		14'b10000000011010:	sigmoid = 21'b000000000000000000001;
		14'b10000000011011:	sigmoid = 21'b000000000000000000001;
		14'b10000000011100:	sigmoid = 21'b000000000000000000001;
		14'b10000000011101:	sigmoid = 21'b000000000000000000001;
		14'b10000000011110:	sigmoid = 21'b000000000000000000001;
		14'b10000000011111:	sigmoid = 21'b000000000000000000001;
		14'b10000000100000:	sigmoid = 21'b000000000000000000001;
		14'b10000000100001:	sigmoid = 21'b000000000000000000001;
		14'b10000000100010:	sigmoid = 21'b000000000000000000001;
		14'b10000000100011:	sigmoid = 21'b000000000000000000001;
		14'b10000000100100:	sigmoid = 21'b000000000000000000001;
		14'b10000000100101:	sigmoid = 21'b000000000000000000001;
		14'b10000000100110:	sigmoid = 21'b000000000000000000001;
		14'b10000000100111:	sigmoid = 21'b000000000000000000001;
		14'b10000000101000:	sigmoid = 21'b000000000000000000001;
		14'b10000000101001:	sigmoid = 21'b000000000000000000001;
		14'b10000000101010:	sigmoid = 21'b000000000000000000001;
		14'b10000000101011:	sigmoid = 21'b000000000000000000001;
		14'b10000000101100:	sigmoid = 21'b000000000000000000001;
		14'b10000000101101:	sigmoid = 21'b000000000000000000001;
		14'b10000000101110:	sigmoid = 21'b000000000000000000001;
		14'b10000000101111:	sigmoid = 21'b000000000000000000001;
		14'b10000000110000:	sigmoid = 21'b000000000000000000001;
		14'b10000000110001:	sigmoid = 21'b000000000000000000001;
		14'b10000000110010:	sigmoid = 21'b000000000000000000001;
		14'b10000000110011:	sigmoid = 21'b000000000000000000001;
		14'b10000000110100:	sigmoid = 21'b000000000000000000001;
		14'b10000000110101:	sigmoid = 21'b000000000000000000001;
		14'b10000000110110:	sigmoid = 21'b000000000000000000001;
		14'b10000000110111:	sigmoid = 21'b000000000000000000001;
		14'b10000000111000:	sigmoid = 21'b000000000000000000001;
		14'b10000000111001:	sigmoid = 21'b000000000000000000001;
		14'b10000000111010:	sigmoid = 21'b000000000000000000001;
		14'b10000000111011:	sigmoid = 21'b000000000000000000001;
		14'b10000000111100:	sigmoid = 21'b000000000000000000001;
		14'b10000000111101:	sigmoid = 21'b000000000000000000001;
		14'b10000000111110:	sigmoid = 21'b000000000000000000001;
		14'b10000000111111:	sigmoid = 21'b000000000000000000001;
		14'b10000001000000:	sigmoid = 21'b000000000000000000001;
		14'b10000001000001:	sigmoid = 21'b000000000000000000001;
		14'b10000001000010:	sigmoid = 21'b000000000000000000001;
		14'b10000001000011:	sigmoid = 21'b000000000000000000001;
		14'b10000001000100:	sigmoid = 21'b000000000000000000001;
		14'b10000001000101:	sigmoid = 21'b000000000000000000001;
		14'b10000001000110:	sigmoid = 21'b000000000000000000001;
		14'b10000001000111:	sigmoid = 21'b000000000000000000001;
		14'b10000001001000:	sigmoid = 21'b000000000000000000001;
		14'b10000001001001:	sigmoid = 21'b000000000000000000001;
		14'b10000001001010:	sigmoid = 21'b000000000000000000001;
		14'b10000001001011:	sigmoid = 21'b000000000000000000001;
		14'b10000001001100:	sigmoid = 21'b000000000000000000001;
		14'b10000001001101:	sigmoid = 21'b000000000000000000001;
		14'b10000001001110:	sigmoid = 21'b000000000000000000001;
		14'b10000001001111:	sigmoid = 21'b000000000000000000001;
		14'b10000001010000:	sigmoid = 21'b000000000000000000001;
		14'b10000001010001:	sigmoid = 21'b000000000000000000001;
		14'b10000001010010:	sigmoid = 21'b000000000000000000001;
		14'b10000001010011:	sigmoid = 21'b000000000000000000001;
		14'b10000001010100:	sigmoid = 21'b000000000000000000001;
		14'b10000001010101:	sigmoid = 21'b000000000000000000001;
		14'b10000001010110:	sigmoid = 21'b000000000000000000001;
		14'b10000001010111:	sigmoid = 21'b000000000000000000001;
		14'b10000001011000:	sigmoid = 21'b000000000000000000001;
		14'b10000001011001:	sigmoid = 21'b000000000000000000001;
		14'b10000001011010:	sigmoid = 21'b000000000000000000001;
		14'b10000001011011:	sigmoid = 21'b000000000000000000001;
		14'b10000001011100:	sigmoid = 21'b000000000000000000001;
		14'b10000001011101:	sigmoid = 21'b000000000000000000001;
		14'b10000001011110:	sigmoid = 21'b000000000000000000001;
		14'b10000001011111:	sigmoid = 21'b000000000000000000001;
		14'b10000001100000:	sigmoid = 21'b000000000000000000001;
		14'b10000001100001:	sigmoid = 21'b000000000000000000001;
		14'b10000001100010:	sigmoid = 21'b000000000000000000001;
		14'b10000001100011:	sigmoid = 21'b000000000000000000001;
		14'b10000001100100:	sigmoid = 21'b000000000000000000001;
		14'b10000001100101:	sigmoid = 21'b000000000000000000001;
		14'b10000001100110:	sigmoid = 21'b000000000000000000001;
		14'b10000001100111:	sigmoid = 21'b000000000000000000001;
		14'b10000001101000:	sigmoid = 21'b000000000000000000001;
		14'b10000001101001:	sigmoid = 21'b000000000000000000001;
		14'b10000001101010:	sigmoid = 21'b000000000000000000001;
		14'b10000001101011:	sigmoid = 21'b000000000000000000001;
		14'b10000001101100:	sigmoid = 21'b000000000000000000001;
		14'b10000001101101:	sigmoid = 21'b000000000000000000001;
		14'b10000001101110:	sigmoid = 21'b000000000000000000001;
		14'b10000001101111:	sigmoid = 21'b000000000000000000001;
		14'b10000001110000:	sigmoid = 21'b000000000000000000001;
		14'b10000001110001:	sigmoid = 21'b000000000000000000001;
		14'b10000001110010:	sigmoid = 21'b000000000000000000001;
		14'b10000001110011:	sigmoid = 21'b000000000000000000001;
		14'b10000001110100:	sigmoid = 21'b000000000000000000001;
		14'b10000001110101:	sigmoid = 21'b000000000000000000001;
		14'b10000001110110:	sigmoid = 21'b000000000000000000001;
		14'b10000001110111:	sigmoid = 21'b000000000000000000001;
		14'b10000001111000:	sigmoid = 21'b000000000000000000001;
		14'b10000001111001:	sigmoid = 21'b000000000000000000001;
		14'b10000001111010:	sigmoid = 21'b000000000000000000001;
		14'b10000001111011:	sigmoid = 21'b000000000000000000001;
		14'b10000001111100:	sigmoid = 21'b000000000000000000001;
		14'b10000001111101:	sigmoid = 21'b000000000000000000001;
		14'b10000001111110:	sigmoid = 21'b000000000000000000001;
		14'b10000001111111:	sigmoid = 21'b000000000000000000001;
		14'b10000010000000:	sigmoid = 21'b000000000000000000001;
		14'b10000010000001:	sigmoid = 21'b000000000000000000001;
		14'b10000010000010:	sigmoid = 21'b000000000000000000001;
		14'b10000010000011:	sigmoid = 21'b000000000000000000001;
		14'b10000010000100:	sigmoid = 21'b000000000000000000001;
		14'b10000010000101:	sigmoid = 21'b000000000000000000001;
		14'b10000010000110:	sigmoid = 21'b000000000000000000001;
		14'b10000010000111:	sigmoid = 21'b000000000000000000001;
		14'b10000010001000:	sigmoid = 21'b000000000000000000001;
		14'b10000010001001:	sigmoid = 21'b000000000000000000001;
		14'b10000010001010:	sigmoid = 21'b000000000000000000001;
		14'b10000010001011:	sigmoid = 21'b000000000000000000001;
		14'b10000010001100:	sigmoid = 21'b000000000000000000001;
		14'b10000010001101:	sigmoid = 21'b000000000000000000001;
		14'b10000010001110:	sigmoid = 21'b000000000000000000001;
		14'b10000010001111:	sigmoid = 21'b000000000000000000001;
		14'b10000010010000:	sigmoid = 21'b000000000000000000001;
		14'b10000010010001:	sigmoid = 21'b000000000000000000001;
		14'b10000010010010:	sigmoid = 21'b000000000000000000001;
		14'b10000010010011:	sigmoid = 21'b000000000000000000001;
		14'b10000010010100:	sigmoid = 21'b000000000000000000001;
		14'b10000010010101:	sigmoid = 21'b000000000000000000001;
		14'b10000010010110:	sigmoid = 21'b000000000000000000001;
		14'b10000010010111:	sigmoid = 21'b000000000000000000001;
		14'b10000010011000:	sigmoid = 21'b000000000000000000001;
		14'b10000010011001:	sigmoid = 21'b000000000000000000001;
		14'b10000010011010:	sigmoid = 21'b000000000000000000001;
		14'b10000010011011:	sigmoid = 21'b000000000000000000001;
		14'b10000010011100:	sigmoid = 21'b000000000000000000001;
		14'b10000010011101:	sigmoid = 21'b000000000000000000001;
		14'b10000010011110:	sigmoid = 21'b000000000000000000001;
		14'b10000010011111:	sigmoid = 21'b000000000000000000001;
		14'b10000010100000:	sigmoid = 21'b000000000000000000001;
		14'b10000010100001:	sigmoid = 21'b000000000000000000001;
		14'b10000010100010:	sigmoid = 21'b000000000000000000001;
		14'b10000010100011:	sigmoid = 21'b000000000000000000001;
		14'b10000010100100:	sigmoid = 21'b000000000000000000001;
		14'b10000010100101:	sigmoid = 21'b000000000000000000001;
		14'b10000010100110:	sigmoid = 21'b000000000000000000001;
		14'b10000010100111:	sigmoid = 21'b000000000000000000001;
		14'b10000010101000:	sigmoid = 21'b000000000000000000001;
		14'b10000010101001:	sigmoid = 21'b000000000000000000001;
		14'b10000010101010:	sigmoid = 21'b000000000000000000001;
		14'b10000010101011:	sigmoid = 21'b000000000000000000001;
		14'b10000010101100:	sigmoid = 21'b000000000000000000001;
		14'b10000010101101:	sigmoid = 21'b000000000000000000001;
		14'b10000010101110:	sigmoid = 21'b000000000000000000001;
		14'b10000010101111:	sigmoid = 21'b000000000000000000001;
		14'b10000010110000:	sigmoid = 21'b000000000000000000001;
		14'b10000010110001:	sigmoid = 21'b000000000000000000001;
		14'b10000010110010:	sigmoid = 21'b000000000000000000001;
		14'b10000010110011:	sigmoid = 21'b000000000000000000001;
		14'b10000010110100:	sigmoid = 21'b000000000000000000001;
		14'b10000010110101:	sigmoid = 21'b000000000000000000001;
		14'b10000010110110:	sigmoid = 21'b000000000000000000001;
		14'b10000010110111:	sigmoid = 21'b000000000000000000001;
		14'b10000010111000:	sigmoid = 21'b000000000000000000001;
		14'b10000010111001:	sigmoid = 21'b000000000000000000001;
		14'b10000010111010:	sigmoid = 21'b000000000000000000001;
		14'b10000010111011:	sigmoid = 21'b000000000000000000001;
		14'b10000010111100:	sigmoid = 21'b000000000000000000001;
		14'b10000010111101:	sigmoid = 21'b000000000000000000001;
		14'b10000010111110:	sigmoid = 21'b000000000000000000001;
		14'b10000010111111:	sigmoid = 21'b000000000000000000001;
		14'b10000011000000:	sigmoid = 21'b000000000000000000001;
		14'b10000011000001:	sigmoid = 21'b000000000000000000001;
		14'b10000011000010:	sigmoid = 21'b000000000000000000001;
		14'b10000011000011:	sigmoid = 21'b000000000000000000001;
		14'b10000011000100:	sigmoid = 21'b000000000000000000001;
		14'b10000011000101:	sigmoid = 21'b000000000000000000001;
		14'b10000011000110:	sigmoid = 21'b000000000000000000001;
		14'b10000011000111:	sigmoid = 21'b000000000000000000001;
		14'b10000011001000:	sigmoid = 21'b000000000000000000001;
		14'b10000011001001:	sigmoid = 21'b000000000000000000001;
		14'b10000011001010:	sigmoid = 21'b000000000000000000001;
		14'b10000011001011:	sigmoid = 21'b000000000000000000001;
		14'b10000011001100:	sigmoid = 21'b000000000000000000001;
		14'b10000011001101:	sigmoid = 21'b000000000000000000001;
		14'b10000011001110:	sigmoid = 21'b000000000000000000001;
		14'b10000011001111:	sigmoid = 21'b000000000000000000001;
		14'b10000011010000:	sigmoid = 21'b000000000000000000001;
		14'b10000011010001:	sigmoid = 21'b000000000000000000001;
		14'b10000011010010:	sigmoid = 21'b000000000000000000001;
		14'b10000011010011:	sigmoid = 21'b000000000000000000001;
		14'b10000011010100:	sigmoid = 21'b000000000000000000001;
		14'b10000011010101:	sigmoid = 21'b000000000000000000001;
		14'b10000011010110:	sigmoid = 21'b000000000000000000001;
		14'b10000011010111:	sigmoid = 21'b000000000000000000001;
		14'b10000011011000:	sigmoid = 21'b000000000000000000001;
		14'b10000011011001:	sigmoid = 21'b000000000000000000001;
		14'b10000011011010:	sigmoid = 21'b000000000000000000001;
		14'b10000011011011:	sigmoid = 21'b000000000000000000001;
		14'b10000011011100:	sigmoid = 21'b000000000000000000001;
		14'b10000011011101:	sigmoid = 21'b000000000000000000001;
		14'b10000011011110:	sigmoid = 21'b000000000000000000001;
		14'b10000011011111:	sigmoid = 21'b000000000000000000001;
		14'b10000011100000:	sigmoid = 21'b000000000000000000001;
		14'b10000011100001:	sigmoid = 21'b000000000000000000001;
		14'b10000011100010:	sigmoid = 21'b000000000000000000001;
		14'b10000011100011:	sigmoid = 21'b000000000000000000001;
		14'b10000011100100:	sigmoid = 21'b000000000000000000001;
		14'b10000011100101:	sigmoid = 21'b000000000000000000001;
		14'b10000011100110:	sigmoid = 21'b000000000000000000001;
		14'b10000011100111:	sigmoid = 21'b000000000000000000001;
		14'b10000011101000:	sigmoid = 21'b000000000000000000001;
		14'b10000011101001:	sigmoid = 21'b000000000000000000001;
		14'b10000011101010:	sigmoid = 21'b000000000000000000001;
		14'b10000011101011:	sigmoid = 21'b000000000000000000001;
		14'b10000011101100:	sigmoid = 21'b000000000000000000001;
		14'b10000011101101:	sigmoid = 21'b000000000000000000001;
		14'b10000011101110:	sigmoid = 21'b000000000000000000001;
		14'b10000011101111:	sigmoid = 21'b000000000000000000001;
		14'b10000011110000:	sigmoid = 21'b000000000000000000001;
		14'b10000011110001:	sigmoid = 21'b000000000000000000001;
		14'b10000011110010:	sigmoid = 21'b000000000000000000001;
		14'b10000011110011:	sigmoid = 21'b000000000000000000001;
		14'b10000011110100:	sigmoid = 21'b000000000000000000001;
		14'b10000011110101:	sigmoid = 21'b000000000000000000001;
		14'b10000011110110:	sigmoid = 21'b000000000000000000001;
		14'b10000011110111:	sigmoid = 21'b000000000000000000001;
		14'b10000011111000:	sigmoid = 21'b000000000000000000001;
		14'b10000011111001:	sigmoid = 21'b000000000000000000001;
		14'b10000011111010:	sigmoid = 21'b000000000000000000001;
		14'b10000011111011:	sigmoid = 21'b000000000000000000001;
		14'b10000011111100:	sigmoid = 21'b000000000000000000001;
		14'b10000011111101:	sigmoid = 21'b000000000000000000001;
		14'b10000011111110:	sigmoid = 21'b000000000000000000001;
		14'b10000011111111:	sigmoid = 21'b000000000000000000001;
		14'b10000100000000:	sigmoid = 21'b000000000000000000001;
		14'b10000100000001:	sigmoid = 21'b000000000000000000001;
		14'b10000100000010:	sigmoid = 21'b000000000000000000001;
		14'b10000100000011:	sigmoid = 21'b000000000000000000001;
		14'b10000100000100:	sigmoid = 21'b000000000000000000001;
		14'b10000100000101:	sigmoid = 21'b000000000000000000001;
		14'b10000100000110:	sigmoid = 21'b000000000000000000001;
		14'b10000100000111:	sigmoid = 21'b000000000000000000001;
		14'b10000100001000:	sigmoid = 21'b000000000000000000001;
		14'b10000100001001:	sigmoid = 21'b000000000000000000001;
		14'b10000100001010:	sigmoid = 21'b000000000000000000001;
		14'b10000100001011:	sigmoid = 21'b000000000000000000001;
		14'b10000100001100:	sigmoid = 21'b000000000000000000001;
		14'b10000100001101:	sigmoid = 21'b000000000000000000001;
		14'b10000100001110:	sigmoid = 21'b000000000000000000001;
		14'b10000100001111:	sigmoid = 21'b000000000000000000001;
		14'b10000100010000:	sigmoid = 21'b000000000000000000001;
		14'b10000100010001:	sigmoid = 21'b000000000000000000001;
		14'b10000100010010:	sigmoid = 21'b000000000000000000001;
		14'b10000100010011:	sigmoid = 21'b000000000000000000001;
		14'b10000100010100:	sigmoid = 21'b000000000000000000001;
		14'b10000100010101:	sigmoid = 21'b000000000000000000001;
		14'b10000100010110:	sigmoid = 21'b000000000000000000001;
		14'b10000100010111:	sigmoid = 21'b000000000000000000001;
		14'b10000100011000:	sigmoid = 21'b000000000000000000001;
		14'b10000100011001:	sigmoid = 21'b000000000000000000001;
		14'b10000100011010:	sigmoid = 21'b000000000000000000001;
		14'b10000100011011:	sigmoid = 21'b000000000000000000001;
		14'b10000100011100:	sigmoid = 21'b000000000000000000001;
		14'b10000100011101:	sigmoid = 21'b000000000000000000001;
		14'b10000100011110:	sigmoid = 21'b000000000000000000001;
		14'b10000100011111:	sigmoid = 21'b000000000000000000001;
		14'b10000100100000:	sigmoid = 21'b000000000000000000001;
		14'b10000100100001:	sigmoid = 21'b000000000000000000001;
		14'b10000100100010:	sigmoid = 21'b000000000000000000001;
		14'b10000100100011:	sigmoid = 21'b000000000000000000001;
		14'b10000100100100:	sigmoid = 21'b000000000000000000001;
		14'b10000100100101:	sigmoid = 21'b000000000000000000001;
		14'b10000100100110:	sigmoid = 21'b000000000000000000001;
		14'b10000100100111:	sigmoid = 21'b000000000000000000001;
		14'b10000100101000:	sigmoid = 21'b000000000000000000001;
		14'b10000100101001:	sigmoid = 21'b000000000000000000001;
		14'b10000100101010:	sigmoid = 21'b000000000000000000001;
		14'b10000100101011:	sigmoid = 21'b000000000000000000001;
		14'b10000100101100:	sigmoid = 21'b000000000000000000001;
		14'b10000100101101:	sigmoid = 21'b000000000000000000001;
		14'b10000100101110:	sigmoid = 21'b000000000000000000001;
		14'b10000100101111:	sigmoid = 21'b000000000000000000001;
		14'b10000100110000:	sigmoid = 21'b000000000000000000001;
		14'b10000100110001:	sigmoid = 21'b000000000000000000001;
		14'b10000100110010:	sigmoid = 21'b000000000000000000001;
		14'b10000100110011:	sigmoid = 21'b000000000000000000001;
		14'b10000100110100:	sigmoid = 21'b000000000000000000001;
		14'b10000100110101:	sigmoid = 21'b000000000000000000001;
		14'b10000100110110:	sigmoid = 21'b000000000000000000001;
		14'b10000100110111:	sigmoid = 21'b000000000000000000001;
		14'b10000100111000:	sigmoid = 21'b000000000000000000001;
		14'b10000100111001:	sigmoid = 21'b000000000000000000001;
		14'b10000100111010:	sigmoid = 21'b000000000000000000001;
		14'b10000100111011:	sigmoid = 21'b000000000000000000001;
		14'b10000100111100:	sigmoid = 21'b000000000000000000001;
		14'b10000100111101:	sigmoid = 21'b000000000000000000001;
		14'b10000100111110:	sigmoid = 21'b000000000000000000001;
		14'b10000100111111:	sigmoid = 21'b000000000000000000001;
		14'b10000101000000:	sigmoid = 21'b000000000000000000001;
		14'b10000101000001:	sigmoid = 21'b000000000000000000001;
		14'b10000101000010:	sigmoid = 21'b000000000000000000001;
		14'b10000101000011:	sigmoid = 21'b000000000000000000001;
		14'b10000101000100:	sigmoid = 21'b000000000000000000001;
		14'b10000101000101:	sigmoid = 21'b000000000000000000001;
		14'b10000101000110:	sigmoid = 21'b000000000000000000001;
		14'b10000101000111:	sigmoid = 21'b000000000000000000001;
		14'b10000101001000:	sigmoid = 21'b000000000000000000001;
		14'b10000101001001:	sigmoid = 21'b000000000000000000001;
		14'b10000101001010:	sigmoid = 21'b000000000000000000001;
		14'b10000101001011:	sigmoid = 21'b000000000000000000001;
		14'b10000101001100:	sigmoid = 21'b000000000000000000001;
		14'b10000101001101:	sigmoid = 21'b000000000000000000001;
		14'b10000101001110:	sigmoid = 21'b000000000000000000001;
		14'b10000101001111:	sigmoid = 21'b000000000000000000001;
		14'b10000101010000:	sigmoid = 21'b000000000000000000001;
		14'b10000101010001:	sigmoid = 21'b000000000000000000001;
		14'b10000101010010:	sigmoid = 21'b000000000000000000001;
		14'b10000101010011:	sigmoid = 21'b000000000000000000001;
		14'b10000101010100:	sigmoid = 21'b000000000000000000001;
		14'b10000101010101:	sigmoid = 21'b000000000000000000001;
		14'b10000101010110:	sigmoid = 21'b000000000000000000001;
		14'b10000101010111:	sigmoid = 21'b000000000000000000001;
		14'b10000101011000:	sigmoid = 21'b000000000000000000001;
		14'b10000101011001:	sigmoid = 21'b000000000000000000001;
		14'b10000101011010:	sigmoid = 21'b000000000000000000001;
		14'b10000101011011:	sigmoid = 21'b000000000000000000001;
		14'b10000101011100:	sigmoid = 21'b000000000000000000001;
		14'b10000101011101:	sigmoid = 21'b000000000000000000001;
		14'b10000101011110:	sigmoid = 21'b000000000000000000001;
		14'b10000101011111:	sigmoid = 21'b000000000000000000001;
		14'b10000101100000:	sigmoid = 21'b000000000000000000001;
		14'b10000101100001:	sigmoid = 21'b000000000000000000001;
		14'b10000101100010:	sigmoid = 21'b000000000000000000001;
		14'b10000101100011:	sigmoid = 21'b000000000000000000001;
		14'b10000101100100:	sigmoid = 21'b000000000000000000001;
		14'b10000101100101:	sigmoid = 21'b000000000000000000001;
		14'b10000101100110:	sigmoid = 21'b000000000000000000001;
		14'b10000101100111:	sigmoid = 21'b000000000000000000001;
		14'b10000101101000:	sigmoid = 21'b000000000000000000001;
		14'b10000101101001:	sigmoid = 21'b000000000000000000001;
		14'b10000101101010:	sigmoid = 21'b000000000000000000001;
		14'b10000101101011:	sigmoid = 21'b000000000000000000001;
		14'b10000101101100:	sigmoid = 21'b000000000000000000001;
		14'b10000101101101:	sigmoid = 21'b000000000000000000001;
		14'b10000101101110:	sigmoid = 21'b000000000000000000001;
		14'b10000101101111:	sigmoid = 21'b000000000000000000001;
		14'b10000101110000:	sigmoid = 21'b000000000000000000001;
		14'b10000101110001:	sigmoid = 21'b000000000000000000001;
		14'b10000101110010:	sigmoid = 21'b000000000000000000001;
		14'b10000101110011:	sigmoid = 21'b000000000000000000001;
		14'b10000101110100:	sigmoid = 21'b000000000000000000001;
		14'b10000101110101:	sigmoid = 21'b000000000000000000001;
		14'b10000101110110:	sigmoid = 21'b000000000000000000001;
		14'b10000101110111:	sigmoid = 21'b000000000000000000001;
		14'b10000101111000:	sigmoid = 21'b000000000000000000001;
		14'b10000101111001:	sigmoid = 21'b000000000000000000001;
		14'b10000101111010:	sigmoid = 21'b000000000000000000001;
		14'b10000101111011:	sigmoid = 21'b000000000000000000001;
		14'b10000101111100:	sigmoid = 21'b000000000000000000001;
		14'b10000101111101:	sigmoid = 21'b000000000000000000001;
		14'b10000101111110:	sigmoid = 21'b000000000000000000001;
		14'b10000101111111:	sigmoid = 21'b000000000000000000001;
		14'b10000110000000:	sigmoid = 21'b000000000000000000001;
		14'b10000110000001:	sigmoid = 21'b000000000000000000001;
		14'b10000110000010:	sigmoid = 21'b000000000000000000001;
		14'b10000110000011:	sigmoid = 21'b000000000000000000001;
		14'b10000110000100:	sigmoid = 21'b000000000000000000001;
		14'b10000110000101:	sigmoid = 21'b000000000000000000001;
		14'b10000110000110:	sigmoid = 21'b000000000000000000001;
		14'b10000110000111:	sigmoid = 21'b000000000000000000001;
		14'b10000110001000:	sigmoid = 21'b000000000000000000001;
		14'b10000110001001:	sigmoid = 21'b000000000000000000001;
		14'b10000110001010:	sigmoid = 21'b000000000000000000001;
		14'b10000110001011:	sigmoid = 21'b000000000000000000001;
		14'b10000110001100:	sigmoid = 21'b000000000000000000001;
		14'b10000110001101:	sigmoid = 21'b000000000000000000001;
		14'b10000110001110:	sigmoid = 21'b000000000000000000001;
		14'b10000110001111:	sigmoid = 21'b000000000000000000001;
		14'b10000110010000:	sigmoid = 21'b000000000000000000001;
		14'b10000110010001:	sigmoid = 21'b000000000000000000001;
		14'b10000110010010:	sigmoid = 21'b000000000000000000001;
		14'b10000110010011:	sigmoid = 21'b000000000000000000001;
		14'b10000110010100:	sigmoid = 21'b000000000000000000001;
		14'b10000110010101:	sigmoid = 21'b000000000000000000001;
		14'b10000110010110:	sigmoid = 21'b000000000000000000001;
		14'b10000110010111:	sigmoid = 21'b000000000000000000001;
		14'b10000110011000:	sigmoid = 21'b000000000000000000001;
		14'b10000110011001:	sigmoid = 21'b000000000000000000001;
		14'b10000110011010:	sigmoid = 21'b000000000000000000001;
		14'b10000110011011:	sigmoid = 21'b000000000000000000001;
		14'b10000110011100:	sigmoid = 21'b000000000000000000001;
		14'b10000110011101:	sigmoid = 21'b000000000000000000001;
		14'b10000110011110:	sigmoid = 21'b000000000000000000001;
		14'b10000110011111:	sigmoid = 21'b000000000000000000001;
		14'b10000110100000:	sigmoid = 21'b000000000000000000001;
		14'b10000110100001:	sigmoid = 21'b000000000000000000001;
		14'b10000110100010:	sigmoid = 21'b000000000000000000001;
		14'b10000110100011:	sigmoid = 21'b000000000000000000001;
		14'b10000110100100:	sigmoid = 21'b000000000000000000001;
		14'b10000110100101:	sigmoid = 21'b000000000000000000001;
		14'b10000110100110:	sigmoid = 21'b000000000000000000001;
		14'b10000110100111:	sigmoid = 21'b000000000000000000001;
		14'b10000110101000:	sigmoid = 21'b000000000000000000001;
		14'b10000110101001:	sigmoid = 21'b000000000000000000001;
		14'b10000110101010:	sigmoid = 21'b000000000000000000001;
		14'b10000110101011:	sigmoid = 21'b000000000000000000001;
		14'b10000110101100:	sigmoid = 21'b000000000000000000001;
		14'b10000110101101:	sigmoid = 21'b000000000000000000001;
		14'b10000110101110:	sigmoid = 21'b000000000000000000001;
		14'b10000110101111:	sigmoid = 21'b000000000000000000001;
		14'b10000110110000:	sigmoid = 21'b000000000000000000001;
		14'b10000110110001:	sigmoid = 21'b000000000000000000001;
		14'b10000110110010:	sigmoid = 21'b000000000000000000001;
		14'b10000110110011:	sigmoid = 21'b000000000000000000001;
		14'b10000110110100:	sigmoid = 21'b000000000000000000001;
		14'b10000110110101:	sigmoid = 21'b000000000000000000001;
		14'b10000110110110:	sigmoid = 21'b000000000000000000001;
		14'b10000110110111:	sigmoid = 21'b000000000000000000001;
		14'b10000110111000:	sigmoid = 21'b000000000000000000001;
		14'b10000110111001:	sigmoid = 21'b000000000000000000001;
		14'b10000110111010:	sigmoid = 21'b000000000000000000001;
		14'b10000110111011:	sigmoid = 21'b000000000000000000001;
		14'b10000110111100:	sigmoid = 21'b000000000000000000001;
		14'b10000110111101:	sigmoid = 21'b000000000000000000001;
		14'b10000110111110:	sigmoid = 21'b000000000000000000001;
		14'b10000110111111:	sigmoid = 21'b000000000000000000001;
		14'b10000111000000:	sigmoid = 21'b000000000000000000001;
		14'b10000111000001:	sigmoid = 21'b000000000000000000001;
		14'b10000111000010:	sigmoid = 21'b000000000000000000001;
		14'b10000111000011:	sigmoid = 21'b000000000000000000001;
		14'b10000111000100:	sigmoid = 21'b000000000000000000001;
		14'b10000111000101:	sigmoid = 21'b000000000000000000001;
		14'b10000111000110:	sigmoid = 21'b000000000000000000001;
		14'b10000111000111:	sigmoid = 21'b000000000000000000001;
		14'b10000111001000:	sigmoid = 21'b000000000000000000001;
		14'b10000111001001:	sigmoid = 21'b000000000000000000001;
		14'b10000111001010:	sigmoid = 21'b000000000000000000001;
		14'b10000111001011:	sigmoid = 21'b000000000000000000001;
		14'b10000111001100:	sigmoid = 21'b000000000000000000001;
		14'b10000111001101:	sigmoid = 21'b000000000000000000001;
		14'b10000111001110:	sigmoid = 21'b000000000000000000001;
		14'b10000111001111:	sigmoid = 21'b000000000000000000001;
		14'b10000111010000:	sigmoid = 21'b000000000000000000001;
		14'b10000111010001:	sigmoid = 21'b000000000000000000001;
		14'b10000111010010:	sigmoid = 21'b000000000000000000001;
		14'b10000111010011:	sigmoid = 21'b000000000000000000001;
		14'b10000111010100:	sigmoid = 21'b000000000000000000001;
		14'b10000111010101:	sigmoid = 21'b000000000000000000001;
		14'b10000111010110:	sigmoid = 21'b000000000000000000001;
		14'b10000111010111:	sigmoid = 21'b000000000000000000001;
		14'b10000111011000:	sigmoid = 21'b000000000000000000001;
		14'b10000111011001:	sigmoid = 21'b000000000000000000001;
		14'b10000111011010:	sigmoid = 21'b000000000000000000001;
		14'b10000111011011:	sigmoid = 21'b000000000000000000001;
		14'b10000111011100:	sigmoid = 21'b000000000000000000001;
		14'b10000111011101:	sigmoid = 21'b000000000000000000001;
		14'b10000111011110:	sigmoid = 21'b000000000000000000001;
		14'b10000111011111:	sigmoid = 21'b000000000000000000001;
		14'b10000111100000:	sigmoid = 21'b000000000000000000001;
		14'b10000111100001:	sigmoid = 21'b000000000000000000001;
		14'b10000111100010:	sigmoid = 21'b000000000000000000001;
		14'b10000111100011:	sigmoid = 21'b000000000000000000001;
		14'b10000111100100:	sigmoid = 21'b000000000000000000001;
		14'b10000111100101:	sigmoid = 21'b000000000000000000001;
		14'b10000111100110:	sigmoid = 21'b000000000000000000001;
		14'b10000111100111:	sigmoid = 21'b000000000000000000001;
		14'b10000111101000:	sigmoid = 21'b000000000000000000001;
		14'b10000111101001:	sigmoid = 21'b000000000000000000001;
		14'b10000111101010:	sigmoid = 21'b000000000000000000001;
		14'b10000111101011:	sigmoid = 21'b000000000000000000001;
		14'b10000111101100:	sigmoid = 21'b000000000000000000001;
		14'b10000111101101:	sigmoid = 21'b000000000000000000001;
		14'b10000111101110:	sigmoid = 21'b000000000000000000001;
		14'b10000111101111:	sigmoid = 21'b000000000000000000001;
		14'b10000111110000:	sigmoid = 21'b000000000000000000001;
		14'b10000111110001:	sigmoid = 21'b000000000000000000001;
		14'b10000111110010:	sigmoid = 21'b000000000000000000001;
		14'b10000111110011:	sigmoid = 21'b000000000000000000001;
		14'b10000111110100:	sigmoid = 21'b000000000000000000001;
		14'b10000111110101:	sigmoid = 21'b000000000000000000001;
		14'b10000111110110:	sigmoid = 21'b000000000000000000001;
		14'b10000111110111:	sigmoid = 21'b000000000000000000001;
		14'b10000111111000:	sigmoid = 21'b000000000000000000001;
		14'b10000111111001:	sigmoid = 21'b000000000000000000001;
		14'b10000111111010:	sigmoid = 21'b000000000000000000001;
		14'b10000111111011:	sigmoid = 21'b000000000000000000001;
		14'b10000111111100:	sigmoid = 21'b000000000000000000001;
		14'b10000111111101:	sigmoid = 21'b000000000000000000001;
		14'b10000111111110:	sigmoid = 21'b000000000000000000001;
		14'b10000111111111:	sigmoid = 21'b000000000000000000001;
		14'b10001000000000:	sigmoid = 21'b000000000000000000001;
		14'b10001000000001:	sigmoid = 21'b000000000000000000001;
		14'b10001000000010:	sigmoid = 21'b000000000000000000001;
		14'b10001000000011:	sigmoid = 21'b000000000000000000001;
		14'b10001000000100:	sigmoid = 21'b000000000000000000001;
		14'b10001000000101:	sigmoid = 21'b000000000000000000001;
		14'b10001000000110:	sigmoid = 21'b000000000000000000001;
		14'b10001000000111:	sigmoid = 21'b000000000000000000001;
		14'b10001000001000:	sigmoid = 21'b000000000000000000001;
		14'b10001000001001:	sigmoid = 21'b000000000000000000001;
		14'b10001000001010:	sigmoid = 21'b000000000000000000001;
		14'b10001000001011:	sigmoid = 21'b000000000000000000001;
		14'b10001000001100:	sigmoid = 21'b000000000000000000001;
		14'b10001000001101:	sigmoid = 21'b000000000000000000001;
		14'b10001000001110:	sigmoid = 21'b000000000000000000001;
		14'b10001000001111:	sigmoid = 21'b000000000000000000001;
		14'b10001000010000:	sigmoid = 21'b000000000000000000001;
		14'b10001000010001:	sigmoid = 21'b000000000000000000001;
		14'b10001000010010:	sigmoid = 21'b000000000000000000001;
		14'b10001000010011:	sigmoid = 21'b000000000000000000001;
		14'b10001000010100:	sigmoid = 21'b000000000000000000001;
		14'b10001000010101:	sigmoid = 21'b000000000000000000001;
		14'b10001000010110:	sigmoid = 21'b000000000000000000001;
		14'b10001000010111:	sigmoid = 21'b000000000000000000001;
		14'b10001000011000:	sigmoid = 21'b000000000000000000001;
		14'b10001000011001:	sigmoid = 21'b000000000000000000001;
		14'b10001000011010:	sigmoid = 21'b000000000000000000001;
		14'b10001000011011:	sigmoid = 21'b000000000000000000001;
		14'b10001000011100:	sigmoid = 21'b000000000000000000001;
		14'b10001000011101:	sigmoid = 21'b000000000000000000001;
		14'b10001000011110:	sigmoid = 21'b000000000000000000001;
		14'b10001000011111:	sigmoid = 21'b000000000000000000001;
		14'b10001000100000:	sigmoid = 21'b000000000000000000001;
		14'b10001000100001:	sigmoid = 21'b000000000000000000001;
		14'b10001000100010:	sigmoid = 21'b000000000000000000001;
		14'b10001000100011:	sigmoid = 21'b000000000000000000001;
		14'b10001000100100:	sigmoid = 21'b000000000000000000001;
		14'b10001000100101:	sigmoid = 21'b000000000000000000001;
		14'b10001000100110:	sigmoid = 21'b000000000000000000001;
		14'b10001000100111:	sigmoid = 21'b000000000000000000001;
		14'b10001000101000:	sigmoid = 21'b000000000000000000001;
		14'b10001000101001:	sigmoid = 21'b000000000000000000001;
		14'b10001000101010:	sigmoid = 21'b000000000000000000001;
		14'b10001000101011:	sigmoid = 21'b000000000000000000001;
		14'b10001000101100:	sigmoid = 21'b000000000000000000001;
		14'b10001000101101:	sigmoid = 21'b000000000000000000001;
		14'b10001000101110:	sigmoid = 21'b000000000000000000001;
		14'b10001000101111:	sigmoid = 21'b000000000000000000001;
		14'b10001000110000:	sigmoid = 21'b000000000000000000001;
		14'b10001000110001:	sigmoid = 21'b000000000000000000001;
		14'b10001000110010:	sigmoid = 21'b000000000000000000001;
		14'b10001000110011:	sigmoid = 21'b000000000000000000001;
		14'b10001000110100:	sigmoid = 21'b000000000000000000001;
		14'b10001000110101:	sigmoid = 21'b000000000000000000001;
		14'b10001000110110:	sigmoid = 21'b000000000000000000001;
		14'b10001000110111:	sigmoid = 21'b000000000000000000001;
		14'b10001000111000:	sigmoid = 21'b000000000000000000001;
		14'b10001000111001:	sigmoid = 21'b000000000000000000001;
		14'b10001000111010:	sigmoid = 21'b000000000000000000001;
		14'b10001000111011:	sigmoid = 21'b000000000000000000001;
		14'b10001000111100:	sigmoid = 21'b000000000000000000001;
		14'b10001000111101:	sigmoid = 21'b000000000000000000001;
		14'b10001000111110:	sigmoid = 21'b000000000000000000001;
		14'b10001000111111:	sigmoid = 21'b000000000000000000001;
		14'b10001001000000:	sigmoid = 21'b000000000000000000001;
		14'b10001001000001:	sigmoid = 21'b000000000000000000001;
		14'b10001001000010:	sigmoid = 21'b000000000000000000001;
		14'b10001001000011:	sigmoid = 21'b000000000000000000001;
		14'b10001001000100:	sigmoid = 21'b000000000000000000001;
		14'b10001001000101:	sigmoid = 21'b000000000000000000001;
		14'b10001001000110:	sigmoid = 21'b000000000000000000001;
		14'b10001001000111:	sigmoid = 21'b000000000000000000001;
		14'b10001001001000:	sigmoid = 21'b000000000000000000001;
		14'b10001001001001:	sigmoid = 21'b000000000000000000001;
		14'b10001001001010:	sigmoid = 21'b000000000000000000001;
		14'b10001001001011:	sigmoid = 21'b000000000000000000001;
		14'b10001001001100:	sigmoid = 21'b000000000000000000001;
		14'b10001001001101:	sigmoid = 21'b000000000000000000001;
		14'b10001001001110:	sigmoid = 21'b000000000000000000001;
		14'b10001001001111:	sigmoid = 21'b000000000000000000001;
		14'b10001001010000:	sigmoid = 21'b000000000000000000001;
		14'b10001001010001:	sigmoid = 21'b000000000000000000001;
		14'b10001001010010:	sigmoid = 21'b000000000000000000001;
		14'b10001001010011:	sigmoid = 21'b000000000000000000001;
		14'b10001001010100:	sigmoid = 21'b000000000000000000001;
		14'b10001001010101:	sigmoid = 21'b000000000000000000001;
		14'b10001001010110:	sigmoid = 21'b000000000000000000001;
		14'b10001001010111:	sigmoid = 21'b000000000000000000001;
		14'b10001001011000:	sigmoid = 21'b000000000000000000001;
		14'b10001001011001:	sigmoid = 21'b000000000000000000001;
		14'b10001001011010:	sigmoid = 21'b000000000000000000001;
		14'b10001001011011:	sigmoid = 21'b000000000000000000001;
		14'b10001001011100:	sigmoid = 21'b000000000000000000001;
		14'b10001001011101:	sigmoid = 21'b000000000000000000001;
		14'b10001001011110:	sigmoid = 21'b000000000000000000001;
		14'b10001001011111:	sigmoid = 21'b000000000000000000001;
		14'b10001001100000:	sigmoid = 21'b000000000000000000001;
		14'b10001001100001:	sigmoid = 21'b000000000000000000001;
		14'b10001001100010:	sigmoid = 21'b000000000000000000001;
		14'b10001001100011:	sigmoid = 21'b000000000000000000001;
		14'b10001001100100:	sigmoid = 21'b000000000000000000001;
		14'b10001001100101:	sigmoid = 21'b000000000000000000001;
		14'b10001001100110:	sigmoid = 21'b000000000000000000001;
		14'b10001001100111:	sigmoid = 21'b000000000000000000001;
		14'b10001001101000:	sigmoid = 21'b000000000000000000001;
		14'b10001001101001:	sigmoid = 21'b000000000000000000001;
		14'b10001001101010:	sigmoid = 21'b000000000000000000001;
		14'b10001001101011:	sigmoid = 21'b000000000000000000001;
		14'b10001001101100:	sigmoid = 21'b000000000000000000001;
		14'b10001001101101:	sigmoid = 21'b000000000000000000001;
		14'b10001001101110:	sigmoid = 21'b000000000000000000001;
		14'b10001001101111:	sigmoid = 21'b000000000000000000001;
		14'b10001001110000:	sigmoid = 21'b000000000000000000001;
		14'b10001001110001:	sigmoid = 21'b000000000000000000001;
		14'b10001001110010:	sigmoid = 21'b000000000000000000001;
		14'b10001001110011:	sigmoid = 21'b000000000000000000001;
		14'b10001001110100:	sigmoid = 21'b000000000000000000001;
		14'b10001001110101:	sigmoid = 21'b000000000000000000001;
		14'b10001001110110:	sigmoid = 21'b000000000000000000001;
		14'b10001001110111:	sigmoid = 21'b000000000000000000001;
		14'b10001001111000:	sigmoid = 21'b000000000000000000001;
		14'b10001001111001:	sigmoid = 21'b000000000000000000001;
		14'b10001001111010:	sigmoid = 21'b000000000000000000001;
		14'b10001001111011:	sigmoid = 21'b000000000000000000001;
		14'b10001001111100:	sigmoid = 21'b000000000000000000001;
		14'b10001001111101:	sigmoid = 21'b000000000000000000001;
		14'b10001001111110:	sigmoid = 21'b000000000000000000001;
		14'b10001001111111:	sigmoid = 21'b000000000000000000001;
		14'b10001010000000:	sigmoid = 21'b000000000000000000001;
		14'b10001010000001:	sigmoid = 21'b000000000000000000001;
		14'b10001010000010:	sigmoid = 21'b000000000000000000001;
		14'b10001010000011:	sigmoid = 21'b000000000000000000001;
		14'b10001010000100:	sigmoid = 21'b000000000000000000001;
		14'b10001010000101:	sigmoid = 21'b000000000000000000001;
		14'b10001010000110:	sigmoid = 21'b000000000000000000001;
		14'b10001010000111:	sigmoid = 21'b000000000000000000001;
		14'b10001010001000:	sigmoid = 21'b000000000000000000001;
		14'b10001010001001:	sigmoid = 21'b000000000000000000001;
		14'b10001010001010:	sigmoid = 21'b000000000000000000001;
		14'b10001010001011:	sigmoid = 21'b000000000000000000001;
		14'b10001010001100:	sigmoid = 21'b000000000000000000001;
		14'b10001010001101:	sigmoid = 21'b000000000000000000001;
		14'b10001010001110:	sigmoid = 21'b000000000000000000001;
		14'b10001010001111:	sigmoid = 21'b000000000000000000001;
		14'b10001010010000:	sigmoid = 21'b000000000000000000001;
		14'b10001010010001:	sigmoid = 21'b000000000000000000001;
		14'b10001010010010:	sigmoid = 21'b000000000000000000001;
		14'b10001010010011:	sigmoid = 21'b000000000000000000001;
		14'b10001010010100:	sigmoid = 21'b000000000000000000001;
		14'b10001010010101:	sigmoid = 21'b000000000000000000001;
		14'b10001010010110:	sigmoid = 21'b000000000000000000001;
		14'b10001010010111:	sigmoid = 21'b000000000000000000001;
		14'b10001010011000:	sigmoid = 21'b000000000000000000001;
		14'b10001010011001:	sigmoid = 21'b000000000000000000001;
		14'b10001010011010:	sigmoid = 21'b000000000000000000001;
		14'b10001010011011:	sigmoid = 21'b000000000000000000001;
		14'b10001010011100:	sigmoid = 21'b000000000000000000001;
		14'b10001010011101:	sigmoid = 21'b000000000000000000001;
		14'b10001010011110:	sigmoid = 21'b000000000000000000001;
		14'b10001010011111:	sigmoid = 21'b000000000000000000001;
		14'b10001010100000:	sigmoid = 21'b000000000000000000001;
		14'b10001010100001:	sigmoid = 21'b000000000000000000001;
		14'b10001010100010:	sigmoid = 21'b000000000000000000001;
		14'b10001010100011:	sigmoid = 21'b000000000000000000001;
		14'b10001010100100:	sigmoid = 21'b000000000000000000001;
		14'b10001010100101:	sigmoid = 21'b000000000000000000001;
		14'b10001010100110:	sigmoid = 21'b000000000000000000001;
		14'b10001010100111:	sigmoid = 21'b000000000000000000001;
		14'b10001010101000:	sigmoid = 21'b000000000000000000001;
		14'b10001010101001:	sigmoid = 21'b000000000000000000001;
		14'b10001010101010:	sigmoid = 21'b000000000000000000001;
		14'b10001010101011:	sigmoid = 21'b000000000000000000001;
		14'b10001010101100:	sigmoid = 21'b000000000000000000001;
		14'b10001010101101:	sigmoid = 21'b000000000000000000001;
		14'b10001010101110:	sigmoid = 21'b000000000000000000001;
		14'b10001010101111:	sigmoid = 21'b000000000000000000001;
		14'b10001010110000:	sigmoid = 21'b000000000000000000001;
		14'b10001010110001:	sigmoid = 21'b000000000000000000001;
		14'b10001010110010:	sigmoid = 21'b000000000000000000001;
		14'b10001010110011:	sigmoid = 21'b000000000000000000001;
		14'b10001010110100:	sigmoid = 21'b000000000000000000001;
		14'b10001010110101:	sigmoid = 21'b000000000000000000001;
		14'b10001010110110:	sigmoid = 21'b000000000000000000001;
		14'b10001010110111:	sigmoid = 21'b000000000000000000001;
		14'b10001010111000:	sigmoid = 21'b000000000000000000001;
		14'b10001010111001:	sigmoid = 21'b000000000000000000001;
		14'b10001010111010:	sigmoid = 21'b000000000000000000001;
		14'b10001010111011:	sigmoid = 21'b000000000000000000001;
		14'b10001010111100:	sigmoid = 21'b000000000000000000001;
		14'b10001010111101:	sigmoid = 21'b000000000000000000001;
		14'b10001010111110:	sigmoid = 21'b000000000000000000001;
		14'b10001010111111:	sigmoid = 21'b000000000000000000001;
		14'b10001011000000:	sigmoid = 21'b000000000000000000001;
		14'b10001011000001:	sigmoid = 21'b000000000000000000001;
		14'b10001011000010:	sigmoid = 21'b000000000000000000001;
		14'b10001011000011:	sigmoid = 21'b000000000000000000001;
		14'b10001011000100:	sigmoid = 21'b000000000000000000001;
		14'b10001011000101:	sigmoid = 21'b000000000000000000001;
		14'b10001011000110:	sigmoid = 21'b000000000000000000001;
		14'b10001011000111:	sigmoid = 21'b000000000000000000001;
		14'b10001011001000:	sigmoid = 21'b000000000000000000001;
		14'b10001011001001:	sigmoid = 21'b000000000000000000001;
		14'b10001011001010:	sigmoid = 21'b000000000000000000001;
		14'b10001011001011:	sigmoid = 21'b000000000000000000001;
		14'b10001011001100:	sigmoid = 21'b000000000000000000001;
		14'b10001011001101:	sigmoid = 21'b000000000000000000001;
		14'b10001011001110:	sigmoid = 21'b000000000000000000001;
		14'b10001011001111:	sigmoid = 21'b000000000000000000001;
		14'b10001011010000:	sigmoid = 21'b000000000000000000001;
		14'b10001011010001:	sigmoid = 21'b000000000000000000001;
		14'b10001011010010:	sigmoid = 21'b000000000000000000001;
		14'b10001011010011:	sigmoid = 21'b000000000000000000001;
		14'b10001011010100:	sigmoid = 21'b000000000000000000001;
		14'b10001011010101:	sigmoid = 21'b000000000000000000001;
		14'b10001011010110:	sigmoid = 21'b000000000000000000001;
		14'b10001011010111:	sigmoid = 21'b000000000000000000001;
		14'b10001011011000:	sigmoid = 21'b000000000000000000001;
		14'b10001011011001:	sigmoid = 21'b000000000000000000001;
		14'b10001011011010:	sigmoid = 21'b000000000000000000001;
		14'b10001011011011:	sigmoid = 21'b000000000000000000001;
		14'b10001011011100:	sigmoid = 21'b000000000000000000001;
		14'b10001011011101:	sigmoid = 21'b000000000000000000001;
		14'b10001011011110:	sigmoid = 21'b000000000000000000001;
		14'b10001011011111:	sigmoid = 21'b000000000000000000001;
		14'b10001011100000:	sigmoid = 21'b000000000000000000001;
		14'b10001011100001:	sigmoid = 21'b000000000000000000001;
		14'b10001011100010:	sigmoid = 21'b000000000000000000001;
		14'b10001011100011:	sigmoid = 21'b000000000000000000001;
		14'b10001011100100:	sigmoid = 21'b000000000000000000001;
		14'b10001011100101:	sigmoid = 21'b000000000000000000001;
		14'b10001011100110:	sigmoid = 21'b000000000000000000001;
		14'b10001011100111:	sigmoid = 21'b000000000000000000001;
		14'b10001011101000:	sigmoid = 21'b000000000000000000001;
		14'b10001011101001:	sigmoid = 21'b000000000000000000001;
		14'b10001011101010:	sigmoid = 21'b000000000000000000001;
		14'b10001011101011:	sigmoid = 21'b000000000000000000001;
		14'b10001011101100:	sigmoid = 21'b000000000000000000001;
		14'b10001011101101:	sigmoid = 21'b000000000000000000001;
		14'b10001011101110:	sigmoid = 21'b000000000000000000001;
		14'b10001011101111:	sigmoid = 21'b000000000000000000001;
		14'b10001011110000:	sigmoid = 21'b000000000000000000001;
		14'b10001011110001:	sigmoid = 21'b000000000000000000001;
		14'b10001011110010:	sigmoid = 21'b000000000000000000001;
		14'b10001011110011:	sigmoid = 21'b000000000000000000001;
		14'b10001011110100:	sigmoid = 21'b000000000000000000001;
		14'b10001011110101:	sigmoid = 21'b000000000000000000001;
		14'b10001011110110:	sigmoid = 21'b000000000000000000001;
		14'b10001011110111:	sigmoid = 21'b000000000000000000001;
		14'b10001011111000:	sigmoid = 21'b000000000000000000001;
		14'b10001011111001:	sigmoid = 21'b000000000000000000001;
		14'b10001011111010:	sigmoid = 21'b000000000000000000001;
		14'b10001011111011:	sigmoid = 21'b000000000000000000001;
		14'b10001011111100:	sigmoid = 21'b000000000000000000001;
		14'b10001011111101:	sigmoid = 21'b000000000000000000001;
		14'b10001011111110:	sigmoid = 21'b000000000000000000001;
		14'b10001011111111:	sigmoid = 21'b000000000000000000001;
		14'b10001100000000:	sigmoid = 21'b000000000000000000001;
		14'b10001100000001:	sigmoid = 21'b000000000000000000001;
		14'b10001100000010:	sigmoid = 21'b000000000000000000001;
		14'b10001100000011:	sigmoid = 21'b000000000000000000001;
		14'b10001100000100:	sigmoid = 21'b000000000000000000001;
		14'b10001100000101:	sigmoid = 21'b000000000000000000001;
		14'b10001100000110:	sigmoid = 21'b000000000000000000001;
		14'b10001100000111:	sigmoid = 21'b000000000000000000001;
		14'b10001100001000:	sigmoid = 21'b000000000000000000001;
		14'b10001100001001:	sigmoid = 21'b000000000000000000001;
		14'b10001100001010:	sigmoid = 21'b000000000000000000001;
		14'b10001100001011:	sigmoid = 21'b000000000000000000001;
		14'b10001100001100:	sigmoid = 21'b000000000000000000001;
		14'b10001100001101:	sigmoid = 21'b000000000000000000001;
		14'b10001100001110:	sigmoid = 21'b000000000000000000001;
		14'b10001100001111:	sigmoid = 21'b000000000000000000001;
		14'b10001100010000:	sigmoid = 21'b000000000000000000001;
		14'b10001100010001:	sigmoid = 21'b000000000000000000001;
		14'b10001100010010:	sigmoid = 21'b000000000000000000001;
		14'b10001100010011:	sigmoid = 21'b000000000000000000001;
		14'b10001100010100:	sigmoid = 21'b000000000000000000001;
		14'b10001100010101:	sigmoid = 21'b000000000000000000001;
		14'b10001100010110:	sigmoid = 21'b000000000000000000001;
		14'b10001100010111:	sigmoid = 21'b000000000000000000001;
		14'b10001100011000:	sigmoid = 21'b000000000000000000001;
		14'b10001100011001:	sigmoid = 21'b000000000000000000001;
		14'b10001100011010:	sigmoid = 21'b000000000000000000001;
		14'b10001100011011:	sigmoid = 21'b000000000000000000001;
		14'b10001100011100:	sigmoid = 21'b000000000000000000001;
		14'b10001100011101:	sigmoid = 21'b000000000000000000001;
		14'b10001100011110:	sigmoid = 21'b000000000000000000001;
		14'b10001100011111:	sigmoid = 21'b000000000000000000001;
		14'b10001100100000:	sigmoid = 21'b000000000000000000001;
		14'b10001100100001:	sigmoid = 21'b000000000000000000001;
		14'b10001100100010:	sigmoid = 21'b000000000000000000001;
		14'b10001100100011:	sigmoid = 21'b000000000000000000001;
		14'b10001100100100:	sigmoid = 21'b000000000000000000001;
		14'b10001100100101:	sigmoid = 21'b000000000000000000001;
		14'b10001100100110:	sigmoid = 21'b000000000000000000001;
		14'b10001100100111:	sigmoid = 21'b000000000000000000001;
		14'b10001100101000:	sigmoid = 21'b000000000000000000001;
		14'b10001100101001:	sigmoid = 21'b000000000000000000001;
		14'b10001100101010:	sigmoid = 21'b000000000000000000001;
		14'b10001100101011:	sigmoid = 21'b000000000000000000001;
		14'b10001100101100:	sigmoid = 21'b000000000000000000001;
		14'b10001100101101:	sigmoid = 21'b000000000000000000001;
		14'b10001100101110:	sigmoid = 21'b000000000000000000001;
		14'b10001100101111:	sigmoid = 21'b000000000000000000001;
		14'b10001100110000:	sigmoid = 21'b000000000000000000001;
		14'b10001100110001:	sigmoid = 21'b000000000000000000001;
		14'b10001100110010:	sigmoid = 21'b000000000000000000001;
		14'b10001100110011:	sigmoid = 21'b000000000000000000001;
		14'b10001100110100:	sigmoid = 21'b000000000000000000001;
		14'b10001100110101:	sigmoid = 21'b000000000000000000001;
		14'b10001100110110:	sigmoid = 21'b000000000000000000001;
		14'b10001100110111:	sigmoid = 21'b000000000000000000001;
		14'b10001100111000:	sigmoid = 21'b000000000000000000001;
		14'b10001100111001:	sigmoid = 21'b000000000000000000001;
		14'b10001100111010:	sigmoid = 21'b000000000000000000001;
		14'b10001100111011:	sigmoid = 21'b000000000000000000001;
		14'b10001100111100:	sigmoid = 21'b000000000000000000001;
		14'b10001100111101:	sigmoid = 21'b000000000000000000001;
		14'b10001100111110:	sigmoid = 21'b000000000000000000001;
		14'b10001100111111:	sigmoid = 21'b000000000000000000001;
		14'b10001101000000:	sigmoid = 21'b000000000000000000001;
		14'b10001101000001:	sigmoid = 21'b000000000000000000001;
		14'b10001101000010:	sigmoid = 21'b000000000000000000001;
		14'b10001101000011:	sigmoid = 21'b000000000000000000001;
		14'b10001101000100:	sigmoid = 21'b000000000000000000001;
		14'b10001101000101:	sigmoid = 21'b000000000000000000001;
		14'b10001101000110:	sigmoid = 21'b000000000000000000001;
		14'b10001101000111:	sigmoid = 21'b000000000000000000001;
		14'b10001101001000:	sigmoid = 21'b000000000000000000001;
		14'b10001101001001:	sigmoid = 21'b000000000000000000001;
		14'b10001101001010:	sigmoid = 21'b000000000000000000001;
		14'b10001101001011:	sigmoid = 21'b000000000000000000001;
		14'b10001101001100:	sigmoid = 21'b000000000000000000001;
		14'b10001101001101:	sigmoid = 21'b000000000000000000001;
		14'b10001101001110:	sigmoid = 21'b000000000000000000001;
		14'b10001101001111:	sigmoid = 21'b000000000000000000001;
		14'b10001101010000:	sigmoid = 21'b000000000000000000001;
		14'b10001101010001:	sigmoid = 21'b000000000000000000001;
		14'b10001101010010:	sigmoid = 21'b000000000000000000001;
		14'b10001101010011:	sigmoid = 21'b000000000000000000001;
		14'b10001101010100:	sigmoid = 21'b000000000000000000001;
		14'b10001101010101:	sigmoid = 21'b000000000000000000001;
		14'b10001101010110:	sigmoid = 21'b000000000000000000001;
		14'b10001101010111:	sigmoid = 21'b000000000000000000001;
		14'b10001101011000:	sigmoid = 21'b000000000000000000001;
		14'b10001101011001:	sigmoid = 21'b000000000000000000001;
		14'b10001101011010:	sigmoid = 21'b000000000000000000001;
		14'b10001101011011:	sigmoid = 21'b000000000000000000001;
		14'b10001101011100:	sigmoid = 21'b000000000000000000001;
		14'b10001101011101:	sigmoid = 21'b000000000000000000001;
		14'b10001101011110:	sigmoid = 21'b000000000000000000001;
		14'b10001101011111:	sigmoid = 21'b000000000000000000001;
		14'b10001101100000:	sigmoid = 21'b000000000000000000001;
		14'b10001101100001:	sigmoid = 21'b000000000000000000001;
		14'b10001101100010:	sigmoid = 21'b000000000000000000001;
		14'b10001101100011:	sigmoid = 21'b000000000000000000001;
		14'b10001101100100:	sigmoid = 21'b000000000000000000001;
		14'b10001101100101:	sigmoid = 21'b000000000000000000001;
		14'b10001101100110:	sigmoid = 21'b000000000000000000001;
		14'b10001101100111:	sigmoid = 21'b000000000000000000001;
		14'b10001101101000:	sigmoid = 21'b000000000000000000001;
		14'b10001101101001:	sigmoid = 21'b000000000000000000001;
		14'b10001101101010:	sigmoid = 21'b000000000000000000001;
		14'b10001101101011:	sigmoid = 21'b000000000000000000001;
		14'b10001101101100:	sigmoid = 21'b000000000000000000001;
		14'b10001101101101:	sigmoid = 21'b000000000000000000001;
		14'b10001101101110:	sigmoid = 21'b000000000000000000001;
		14'b10001101101111:	sigmoid = 21'b000000000000000000001;
		14'b10001101110000:	sigmoid = 21'b000000000000000000001;
		14'b10001101110001:	sigmoid = 21'b000000000000000000001;
		14'b10001101110010:	sigmoid = 21'b000000000000000000001;
		14'b10001101110011:	sigmoid = 21'b000000000000000000001;
		14'b10001101110100:	sigmoid = 21'b000000000000000000001;
		14'b10001101110101:	sigmoid = 21'b000000000000000000001;
		14'b10001101110110:	sigmoid = 21'b000000000000000000001;
		14'b10001101110111:	sigmoid = 21'b000000000000000000001;
		14'b10001101111000:	sigmoid = 21'b000000000000000000001;
		14'b10001101111001:	sigmoid = 21'b000000000000000000001;
		14'b10001101111010:	sigmoid = 21'b000000000000000000001;
		14'b10001101111011:	sigmoid = 21'b000000000000000000001;
		14'b10001101111100:	sigmoid = 21'b000000000000000000001;
		14'b10001101111101:	sigmoid = 21'b000000000000000000001;
		14'b10001101111110:	sigmoid = 21'b000000000000000000001;
		14'b10001101111111:	sigmoid = 21'b000000000000000000001;
		14'b10001110000000:	sigmoid = 21'b000000000000000000001;
		14'b10001110000001:	sigmoid = 21'b000000000000000000001;
		14'b10001110000010:	sigmoid = 21'b000000000000000000001;
		14'b10001110000011:	sigmoid = 21'b000000000000000000001;
		14'b10001110000100:	sigmoid = 21'b000000000000000000001;
		14'b10001110000101:	sigmoid = 21'b000000000000000000001;
		14'b10001110000110:	sigmoid = 21'b000000000000000000001;
		14'b10001110000111:	sigmoid = 21'b000000000000000000001;
		14'b10001110001000:	sigmoid = 21'b000000000000000000001;
		14'b10001110001001:	sigmoid = 21'b000000000000000000001;
		14'b10001110001010:	sigmoid = 21'b000000000000000000001;
		14'b10001110001011:	sigmoid = 21'b000000000000000000001;
		14'b10001110001100:	sigmoid = 21'b000000000000000000001;
		14'b10001110001101:	sigmoid = 21'b000000000000000000001;
		14'b10001110001110:	sigmoid = 21'b000000000000000000001;
		14'b10001110001111:	sigmoid = 21'b000000000000000000001;
		14'b10001110010000:	sigmoid = 21'b000000000000000000001;
		14'b10001110010001:	sigmoid = 21'b000000000000000000001;
		14'b10001110010010:	sigmoid = 21'b000000000000000000001;
		14'b10001110010011:	sigmoid = 21'b000000000000000000001;
		14'b10001110010100:	sigmoid = 21'b000000000000000000001;
		14'b10001110010101:	sigmoid = 21'b000000000000000000001;
		14'b10001110010110:	sigmoid = 21'b000000000000000000001;
		14'b10001110010111:	sigmoid = 21'b000000000000000000001;
		14'b10001110011000:	sigmoid = 21'b000000000000000000001;
		14'b10001110011001:	sigmoid = 21'b000000000000000000001;
		14'b10001110011010:	sigmoid = 21'b000000000000000000001;
		14'b10001110011011:	sigmoid = 21'b000000000000000000001;
		14'b10001110011100:	sigmoid = 21'b000000000000000000001;
		14'b10001110011101:	sigmoid = 21'b000000000000000000001;
		14'b10001110011110:	sigmoid = 21'b000000000000000000001;
		14'b10001110011111:	sigmoid = 21'b000000000000000000001;
		14'b10001110100000:	sigmoid = 21'b000000000000000000001;
		14'b10001110100001:	sigmoid = 21'b000000000000000000001;
		14'b10001110100010:	sigmoid = 21'b000000000000000000001;
		14'b10001110100011:	sigmoid = 21'b000000000000000000001;
		14'b10001110100100:	sigmoid = 21'b000000000000000000001;
		14'b10001110100101:	sigmoid = 21'b000000000000000000001;
		14'b10001110100110:	sigmoid = 21'b000000000000000000001;
		14'b10001110100111:	sigmoid = 21'b000000000000000000001;
		14'b10001110101000:	sigmoid = 21'b000000000000000000001;
		14'b10001110101001:	sigmoid = 21'b000000000000000000001;
		14'b10001110101010:	sigmoid = 21'b000000000000000000001;
		14'b10001110101011:	sigmoid = 21'b000000000000000000001;
		14'b10001110101100:	sigmoid = 21'b000000000000000000001;
		14'b10001110101101:	sigmoid = 21'b000000000000000000001;
		14'b10001110101110:	sigmoid = 21'b000000000000000000001;
		14'b10001110101111:	sigmoid = 21'b000000000000000000001;
		14'b10001110110000:	sigmoid = 21'b000000000000000000001;
		14'b10001110110001:	sigmoid = 21'b000000000000000000001;
		14'b10001110110010:	sigmoid = 21'b000000000000000000001;
		14'b10001110110011:	sigmoid = 21'b000000000000000000001;
		14'b10001110110100:	sigmoid = 21'b000000000000000000001;
		14'b10001110110101:	sigmoid = 21'b000000000000000000001;
		14'b10001110110110:	sigmoid = 21'b000000000000000000001;
		14'b10001110110111:	sigmoid = 21'b000000000000000000001;
		14'b10001110111000:	sigmoid = 21'b000000000000000000001;
		14'b10001110111001:	sigmoid = 21'b000000000000000000001;
		14'b10001110111010:	sigmoid = 21'b000000000000000000001;
		14'b10001110111011:	sigmoid = 21'b000000000000000000001;
		14'b10001110111100:	sigmoid = 21'b000000000000000000001;
		14'b10001110111101:	sigmoid = 21'b000000000000000000001;
		14'b10001110111110:	sigmoid = 21'b000000000000000000001;
		14'b10001110111111:	sigmoid = 21'b000000000000000000001;
		14'b10001111000000:	sigmoid = 21'b000000000000000000001;
		14'b10001111000001:	sigmoid = 21'b000000000000000000001;
		14'b10001111000010:	sigmoid = 21'b000000000000000000001;
		14'b10001111000011:	sigmoid = 21'b000000000000000000001;
		14'b10001111000100:	sigmoid = 21'b000000000000000000001;
		14'b10001111000101:	sigmoid = 21'b000000000000000000001;
		14'b10001111000110:	sigmoid = 21'b000000000000000000001;
		14'b10001111000111:	sigmoid = 21'b000000000000000000001;
		14'b10001111001000:	sigmoid = 21'b000000000000000000001;
		14'b10001111001001:	sigmoid = 21'b000000000000000000001;
		14'b10001111001010:	sigmoid = 21'b000000000000000000001;
		14'b10001111001011:	sigmoid = 21'b000000000000000000001;
		14'b10001111001100:	sigmoid = 21'b000000000000000000001;
		14'b10001111001101:	sigmoid = 21'b000000000000000000001;
		14'b10001111001110:	sigmoid = 21'b000000000000000000001;
		14'b10001111001111:	sigmoid = 21'b000000000000000000001;
		14'b10001111010000:	sigmoid = 21'b000000000000000000001;
		14'b10001111010001:	sigmoid = 21'b000000000000000000001;
		14'b10001111010010:	sigmoid = 21'b000000000000000000001;
		14'b10001111010011:	sigmoid = 21'b000000000000000000001;
		14'b10001111010100:	sigmoid = 21'b000000000000000000001;
		14'b10001111010101:	sigmoid = 21'b000000000000000000001;
		14'b10001111010110:	sigmoid = 21'b000000000000000000001;
		14'b10001111010111:	sigmoid = 21'b000000000000000000001;
		14'b10001111011000:	sigmoid = 21'b000000000000000000001;
		14'b10001111011001:	sigmoid = 21'b000000000000000000001;
		14'b10001111011010:	sigmoid = 21'b000000000000000000001;
		14'b10001111011011:	sigmoid = 21'b000000000000000000001;
		14'b10001111011100:	sigmoid = 21'b000000000000000000001;
		14'b10001111011101:	sigmoid = 21'b000000000000000000001;
		14'b10001111011110:	sigmoid = 21'b000000000000000000001;
		14'b10001111011111:	sigmoid = 21'b000000000000000000001;
		14'b10001111100000:	sigmoid = 21'b000000000000000000001;
		14'b10001111100001:	sigmoid = 21'b000000000000000000001;
		14'b10001111100010:	sigmoid = 21'b000000000000000000001;
		14'b10001111100011:	sigmoid = 21'b000000000000000000001;
		14'b10001111100100:	sigmoid = 21'b000000000000000000001;
		14'b10001111100101:	sigmoid = 21'b000000000000000000001;
		14'b10001111100110:	sigmoid = 21'b000000000000000000001;
		14'b10001111100111:	sigmoid = 21'b000000000000000000001;
		14'b10001111101000:	sigmoid = 21'b000000000000000000001;
		14'b10001111101001:	sigmoid = 21'b000000000000000000001;
		14'b10001111101010:	sigmoid = 21'b000000000000000000001;
		14'b10001111101011:	sigmoid = 21'b000000000000000000001;
		14'b10001111101100:	sigmoid = 21'b000000000000000000001;
		14'b10001111101101:	sigmoid = 21'b000000000000000000001;
		14'b10001111101110:	sigmoid = 21'b000000000000000000001;
		14'b10001111101111:	sigmoid = 21'b000000000000000000001;
		14'b10001111110000:	sigmoid = 21'b000000000000000000001;
		14'b10001111110001:	sigmoid = 21'b000000000000000000001;
		14'b10001111110010:	sigmoid = 21'b000000000000000000001;
		14'b10001111110011:	sigmoid = 21'b000000000000000000001;
		14'b10001111110100:	sigmoid = 21'b000000000000000000001;
		14'b10001111110101:	sigmoid = 21'b000000000000000000001;
		14'b10001111110110:	sigmoid = 21'b000000000000000000001;
		14'b10001111110111:	sigmoid = 21'b000000000000000000001;
		14'b10001111111000:	sigmoid = 21'b000000000000000000001;
		14'b10001111111001:	sigmoid = 21'b000000000000000000001;
		14'b10001111111010:	sigmoid = 21'b000000000000000000001;
		14'b10001111111011:	sigmoid = 21'b000000000000000000001;
		14'b10001111111100:	sigmoid = 21'b000000000000000000001;
		14'b10001111111101:	sigmoid = 21'b000000000000000000001;
		14'b10001111111110:	sigmoid = 21'b000000000000000000001;
		14'b10001111111111:	sigmoid = 21'b000000000000000000001;
		14'b10010000000000:	sigmoid = 21'b000000000000000000001;
		14'b10010000000001:	sigmoid = 21'b000000000000000000001;
		14'b10010000000010:	sigmoid = 21'b000000000000000000001;
		14'b10010000000011:	sigmoid = 21'b000000000000000000001;
		14'b10010000000100:	sigmoid = 21'b000000000000000000001;
		14'b10010000000101:	sigmoid = 21'b000000000000000000001;
		14'b10010000000110:	sigmoid = 21'b000000000000000000001;
		14'b10010000000111:	sigmoid = 21'b000000000000000000001;
		14'b10010000001000:	sigmoid = 21'b000000000000000000001;
		14'b10010000001001:	sigmoid = 21'b000000000000000000001;
		14'b10010000001010:	sigmoid = 21'b000000000000000000001;
		14'b10010000001011:	sigmoid = 21'b000000000000000000001;
		14'b10010000001100:	sigmoid = 21'b000000000000000000001;
		14'b10010000001101:	sigmoid = 21'b000000000000000000001;
		14'b10010000001110:	sigmoid = 21'b000000000000000000001;
		14'b10010000001111:	sigmoid = 21'b000000000000000000001;
		14'b10010000010000:	sigmoid = 21'b000000000000000000001;
		14'b10010000010001:	sigmoid = 21'b000000000000000000001;
		14'b10010000010010:	sigmoid = 21'b000000000000000000001;
		14'b10010000010011:	sigmoid = 21'b000000000000000000001;
		14'b10010000010100:	sigmoid = 21'b000000000000000000001;
		14'b10010000010101:	sigmoid = 21'b000000000000000000001;
		14'b10010000010110:	sigmoid = 21'b000000000000000000001;
		14'b10010000010111:	sigmoid = 21'b000000000000000000001;
		14'b10010000011000:	sigmoid = 21'b000000000000000000001;
		14'b10010000011001:	sigmoid = 21'b000000000000000000001;
		14'b10010000011010:	sigmoid = 21'b000000000000000000001;
		14'b10010000011011:	sigmoid = 21'b000000000000000000001;
		14'b10010000011100:	sigmoid = 21'b000000000000000000001;
		14'b10010000011101:	sigmoid = 21'b000000000000000000001;
		14'b10010000011110:	sigmoid = 21'b000000000000000000001;
		14'b10010000011111:	sigmoid = 21'b000000000000000000001;
		14'b10010000100000:	sigmoid = 21'b000000000000000000001;
		14'b10010000100001:	sigmoid = 21'b000000000000000000001;
		14'b10010000100010:	sigmoid = 21'b000000000000000000001;
		14'b10010000100011:	sigmoid = 21'b000000000000000000001;
		14'b10010000100100:	sigmoid = 21'b000000000000000000001;
		14'b10010000100101:	sigmoid = 21'b000000000000000000001;
		14'b10010000100110:	sigmoid = 21'b000000000000000000001;
		14'b10010000100111:	sigmoid = 21'b000000000000000000001;
		14'b10010000101000:	sigmoid = 21'b000000000000000000001;
		14'b10010000101001:	sigmoid = 21'b000000000000000000001;
		14'b10010000101010:	sigmoid = 21'b000000000000000000001;
		14'b10010000101011:	sigmoid = 21'b000000000000000000001;
		14'b10010000101100:	sigmoid = 21'b000000000000000000001;
		14'b10010000101101:	sigmoid = 21'b000000000000000000001;
		14'b10010000101110:	sigmoid = 21'b000000000000000000001;
		14'b10010000101111:	sigmoid = 21'b000000000000000000001;
		14'b10010000110000:	sigmoid = 21'b000000000000000000001;
		14'b10010000110001:	sigmoid = 21'b000000000000000000001;
		14'b10010000110010:	sigmoid = 21'b000000000000000000001;
		14'b10010000110011:	sigmoid = 21'b000000000000000000001;
		14'b10010000110100:	sigmoid = 21'b000000000000000000001;
		14'b10010000110101:	sigmoid = 21'b000000000000000000001;
		14'b10010000110110:	sigmoid = 21'b000000000000000000001;
		14'b10010000110111:	sigmoid = 21'b000000000000000000001;
		14'b10010000111000:	sigmoid = 21'b000000000000000000001;
		14'b10010000111001:	sigmoid = 21'b000000000000000000001;
		14'b10010000111010:	sigmoid = 21'b000000000000000000001;
		14'b10010000111011:	sigmoid = 21'b000000000000000000001;
		14'b10010000111100:	sigmoid = 21'b000000000000000000001;
		14'b10010000111101:	sigmoid = 21'b000000000000000000001;
		14'b10010000111110:	sigmoid = 21'b000000000000000000001;
		14'b10010000111111:	sigmoid = 21'b000000000000000000001;
		14'b10010001000000:	sigmoid = 21'b000000000000000000001;
		14'b10010001000001:	sigmoid = 21'b000000000000000000001;
		14'b10010001000010:	sigmoid = 21'b000000000000000000001;
		14'b10010001000011:	sigmoid = 21'b000000000000000000001;
		14'b10010001000100:	sigmoid = 21'b000000000000000000001;
		14'b10010001000101:	sigmoid = 21'b000000000000000000001;
		14'b10010001000110:	sigmoid = 21'b000000000000000000001;
		14'b10010001000111:	sigmoid = 21'b000000000000000000010;
		14'b10010001001000:	sigmoid = 21'b000000000000000000010;
		14'b10010001001001:	sigmoid = 21'b000000000000000000010;
		14'b10010001001010:	sigmoid = 21'b000000000000000000010;
		14'b10010001001011:	sigmoid = 21'b000000000000000000010;
		14'b10010001001100:	sigmoid = 21'b000000000000000000010;
		14'b10010001001101:	sigmoid = 21'b000000000000000000010;
		14'b10010001001110:	sigmoid = 21'b000000000000000000010;
		14'b10010001001111:	sigmoid = 21'b000000000000000000010;
		14'b10010001010000:	sigmoid = 21'b000000000000000000010;
		14'b10010001010001:	sigmoid = 21'b000000000000000000010;
		14'b10010001010010:	sigmoid = 21'b000000000000000000010;
		14'b10010001010011:	sigmoid = 21'b000000000000000000010;
		14'b10010001010100:	sigmoid = 21'b000000000000000000010;
		14'b10010001010101:	sigmoid = 21'b000000000000000000010;
		14'b10010001010110:	sigmoid = 21'b000000000000000000010;
		14'b10010001010111:	sigmoid = 21'b000000000000000000010;
		14'b10010001011000:	sigmoid = 21'b000000000000000000010;
		14'b10010001011001:	sigmoid = 21'b000000000000000000010;
		14'b10010001011010:	sigmoid = 21'b000000000000000000010;
		14'b10010001011011:	sigmoid = 21'b000000000000000000010;
		14'b10010001011100:	sigmoid = 21'b000000000000000000010;
		14'b10010001011101:	sigmoid = 21'b000000000000000000010;
		14'b10010001011110:	sigmoid = 21'b000000000000000000010;
		14'b10010001011111:	sigmoid = 21'b000000000000000000010;
		14'b10010001100000:	sigmoid = 21'b000000000000000000010;
		14'b10010001100001:	sigmoid = 21'b000000000000000000010;
		14'b10010001100010:	sigmoid = 21'b000000000000000000010;
		14'b10010001100011:	sigmoid = 21'b000000000000000000010;
		14'b10010001100100:	sigmoid = 21'b000000000000000000010;
		14'b10010001100101:	sigmoid = 21'b000000000000000000010;
		14'b10010001100110:	sigmoid = 21'b000000000000000000010;
		14'b10010001100111:	sigmoid = 21'b000000000000000000010;
		14'b10010001101000:	sigmoid = 21'b000000000000000000010;
		14'b10010001101001:	sigmoid = 21'b000000000000000000010;
		14'b10010001101010:	sigmoid = 21'b000000000000000000010;
		14'b10010001101011:	sigmoid = 21'b000000000000000000010;
		14'b10010001101100:	sigmoid = 21'b000000000000000000010;
		14'b10010001101101:	sigmoid = 21'b000000000000000000010;
		14'b10010001101110:	sigmoid = 21'b000000000000000000010;
		14'b10010001101111:	sigmoid = 21'b000000000000000000010;
		14'b10010001110000:	sigmoid = 21'b000000000000000000010;
		14'b10010001110001:	sigmoid = 21'b000000000000000000010;
		14'b10010001110010:	sigmoid = 21'b000000000000000000010;
		14'b10010001110011:	sigmoid = 21'b000000000000000000010;
		14'b10010001110100:	sigmoid = 21'b000000000000000000010;
		14'b10010001110101:	sigmoid = 21'b000000000000000000010;
		14'b10010001110110:	sigmoid = 21'b000000000000000000010;
		14'b10010001110111:	sigmoid = 21'b000000000000000000010;
		14'b10010001111000:	sigmoid = 21'b000000000000000000010;
		14'b10010001111001:	sigmoid = 21'b000000000000000000010;
		14'b10010001111010:	sigmoid = 21'b000000000000000000010;
		14'b10010001111011:	sigmoid = 21'b000000000000000000010;
		14'b10010001111100:	sigmoid = 21'b000000000000000000010;
		14'b10010001111101:	sigmoid = 21'b000000000000000000010;
		14'b10010001111110:	sigmoid = 21'b000000000000000000010;
		14'b10010001111111:	sigmoid = 21'b000000000000000000010;
		14'b10010010000000:	sigmoid = 21'b000000000000000000010;
		14'b10010010000001:	sigmoid = 21'b000000000000000000010;
		14'b10010010000010:	sigmoid = 21'b000000000000000000010;
		14'b10010010000011:	sigmoid = 21'b000000000000000000010;
		14'b10010010000100:	sigmoid = 21'b000000000000000000010;
		14'b10010010000101:	sigmoid = 21'b000000000000000000010;
		14'b10010010000110:	sigmoid = 21'b000000000000000000010;
		14'b10010010000111:	sigmoid = 21'b000000000000000000010;
		14'b10010010001000:	sigmoid = 21'b000000000000000000010;
		14'b10010010001001:	sigmoid = 21'b000000000000000000010;
		14'b10010010001010:	sigmoid = 21'b000000000000000000010;
		14'b10010010001011:	sigmoid = 21'b000000000000000000010;
		14'b10010010001100:	sigmoid = 21'b000000000000000000010;
		14'b10010010001101:	sigmoid = 21'b000000000000000000010;
		14'b10010010001110:	sigmoid = 21'b000000000000000000010;
		14'b10010010001111:	sigmoid = 21'b000000000000000000010;
		14'b10010010010000:	sigmoid = 21'b000000000000000000010;
		14'b10010010010001:	sigmoid = 21'b000000000000000000010;
		14'b10010010010010:	sigmoid = 21'b000000000000000000010;
		14'b10010010010011:	sigmoid = 21'b000000000000000000010;
		14'b10010010010100:	sigmoid = 21'b000000000000000000010;
		14'b10010010010101:	sigmoid = 21'b000000000000000000010;
		14'b10010010010110:	sigmoid = 21'b000000000000000000010;
		14'b10010010010111:	sigmoid = 21'b000000000000000000010;
		14'b10010010011000:	sigmoid = 21'b000000000000000000010;
		14'b10010010011001:	sigmoid = 21'b000000000000000000010;
		14'b10010010011010:	sigmoid = 21'b000000000000000000010;
		14'b10010010011011:	sigmoid = 21'b000000000000000000010;
		14'b10010010011100:	sigmoid = 21'b000000000000000000010;
		14'b10010010011101:	sigmoid = 21'b000000000000000000010;
		14'b10010010011110:	sigmoid = 21'b000000000000000000010;
		14'b10010010011111:	sigmoid = 21'b000000000000000000010;
		14'b10010010100000:	sigmoid = 21'b000000000000000000010;
		14'b10010010100001:	sigmoid = 21'b000000000000000000010;
		14'b10010010100010:	sigmoid = 21'b000000000000000000010;
		14'b10010010100011:	sigmoid = 21'b000000000000000000010;
		14'b10010010100100:	sigmoid = 21'b000000000000000000010;
		14'b10010010100101:	sigmoid = 21'b000000000000000000010;
		14'b10010010100110:	sigmoid = 21'b000000000000000000010;
		14'b10010010100111:	sigmoid = 21'b000000000000000000010;
		14'b10010010101000:	sigmoid = 21'b000000000000000000010;
		14'b10010010101001:	sigmoid = 21'b000000000000000000010;
		14'b10010010101010:	sigmoid = 21'b000000000000000000010;
		14'b10010010101011:	sigmoid = 21'b000000000000000000010;
		14'b10010010101100:	sigmoid = 21'b000000000000000000010;
		14'b10010010101101:	sigmoid = 21'b000000000000000000010;
		14'b10010010101110:	sigmoid = 21'b000000000000000000010;
		14'b10010010101111:	sigmoid = 21'b000000000000000000010;
		14'b10010010110000:	sigmoid = 21'b000000000000000000010;
		14'b10010010110001:	sigmoid = 21'b000000000000000000010;
		14'b10010010110010:	sigmoid = 21'b000000000000000000010;
		14'b10010010110011:	sigmoid = 21'b000000000000000000010;
		14'b10010010110100:	sigmoid = 21'b000000000000000000010;
		14'b10010010110101:	sigmoid = 21'b000000000000000000010;
		14'b10010010110110:	sigmoid = 21'b000000000000000000010;
		14'b10010010110111:	sigmoid = 21'b000000000000000000010;
		14'b10010010111000:	sigmoid = 21'b000000000000000000010;
		14'b10010010111001:	sigmoid = 21'b000000000000000000010;
		14'b10010010111010:	sigmoid = 21'b000000000000000000010;
		14'b10010010111011:	sigmoid = 21'b000000000000000000010;
		14'b10010010111100:	sigmoid = 21'b000000000000000000010;
		14'b10010010111101:	sigmoid = 21'b000000000000000000010;
		14'b10010010111110:	sigmoid = 21'b000000000000000000010;
		14'b10010010111111:	sigmoid = 21'b000000000000000000010;
		14'b10010011000000:	sigmoid = 21'b000000000000000000010;
		14'b10010011000001:	sigmoid = 21'b000000000000000000010;
		14'b10010011000010:	sigmoid = 21'b000000000000000000010;
		14'b10010011000011:	sigmoid = 21'b000000000000000000010;
		14'b10010011000100:	sigmoid = 21'b000000000000000000010;
		14'b10010011000101:	sigmoid = 21'b000000000000000000010;
		14'b10010011000110:	sigmoid = 21'b000000000000000000010;
		14'b10010011000111:	sigmoid = 21'b000000000000000000010;
		14'b10010011001000:	sigmoid = 21'b000000000000000000010;
		14'b10010011001001:	sigmoid = 21'b000000000000000000010;
		14'b10010011001010:	sigmoid = 21'b000000000000000000010;
		14'b10010011001011:	sigmoid = 21'b000000000000000000010;
		14'b10010011001100:	sigmoid = 21'b000000000000000000010;
		14'b10010011001101:	sigmoid = 21'b000000000000000000010;
		14'b10010011001110:	sigmoid = 21'b000000000000000000010;
		14'b10010011001111:	sigmoid = 21'b000000000000000000010;
		14'b10010011010000:	sigmoid = 21'b000000000000000000010;
		14'b10010011010001:	sigmoid = 21'b000000000000000000010;
		14'b10010011010010:	sigmoid = 21'b000000000000000000010;
		14'b10010011010011:	sigmoid = 21'b000000000000000000010;
		14'b10010011010100:	sigmoid = 21'b000000000000000000010;
		14'b10010011010101:	sigmoid = 21'b000000000000000000010;
		14'b10010011010110:	sigmoid = 21'b000000000000000000010;
		14'b10010011010111:	sigmoid = 21'b000000000000000000010;
		14'b10010011011000:	sigmoid = 21'b000000000000000000010;
		14'b10010011011001:	sigmoid = 21'b000000000000000000010;
		14'b10010011011010:	sigmoid = 21'b000000000000000000010;
		14'b10010011011011:	sigmoid = 21'b000000000000000000010;
		14'b10010011011100:	sigmoid = 21'b000000000000000000010;
		14'b10010011011101:	sigmoid = 21'b000000000000000000010;
		14'b10010011011110:	sigmoid = 21'b000000000000000000010;
		14'b10010011011111:	sigmoid = 21'b000000000000000000010;
		14'b10010011100000:	sigmoid = 21'b000000000000000000010;
		14'b10010011100001:	sigmoid = 21'b000000000000000000010;
		14'b10010011100010:	sigmoid = 21'b000000000000000000010;
		14'b10010011100011:	sigmoid = 21'b000000000000000000010;
		14'b10010011100100:	sigmoid = 21'b000000000000000000010;
		14'b10010011100101:	sigmoid = 21'b000000000000000000010;
		14'b10010011100110:	sigmoid = 21'b000000000000000000010;
		14'b10010011100111:	sigmoid = 21'b000000000000000000010;
		14'b10010011101000:	sigmoid = 21'b000000000000000000010;
		14'b10010011101001:	sigmoid = 21'b000000000000000000010;
		14'b10010011101010:	sigmoid = 21'b000000000000000000010;
		14'b10010011101011:	sigmoid = 21'b000000000000000000010;
		14'b10010011101100:	sigmoid = 21'b000000000000000000010;
		14'b10010011101101:	sigmoid = 21'b000000000000000000010;
		14'b10010011101110:	sigmoid = 21'b000000000000000000010;
		14'b10010011101111:	sigmoid = 21'b000000000000000000010;
		14'b10010011110000:	sigmoid = 21'b000000000000000000010;
		14'b10010011110001:	sigmoid = 21'b000000000000000000010;
		14'b10010011110010:	sigmoid = 21'b000000000000000000010;
		14'b10010011110011:	sigmoid = 21'b000000000000000000010;
		14'b10010011110100:	sigmoid = 21'b000000000000000000010;
		14'b10010011110101:	sigmoid = 21'b000000000000000000010;
		14'b10010011110110:	sigmoid = 21'b000000000000000000010;
		14'b10010011110111:	sigmoid = 21'b000000000000000000010;
		14'b10010011111000:	sigmoid = 21'b000000000000000000010;
		14'b10010011111001:	sigmoid = 21'b000000000000000000010;
		14'b10010011111010:	sigmoid = 21'b000000000000000000010;
		14'b10010011111011:	sigmoid = 21'b000000000000000000010;
		14'b10010011111100:	sigmoid = 21'b000000000000000000010;
		14'b10010011111101:	sigmoid = 21'b000000000000000000010;
		14'b10010011111110:	sigmoid = 21'b000000000000000000010;
		14'b10010011111111:	sigmoid = 21'b000000000000000000010;
		14'b10010100000000:	sigmoid = 21'b000000000000000000010;
		14'b10010100000001:	sigmoid = 21'b000000000000000000010;
		14'b10010100000010:	sigmoid = 21'b000000000000000000010;
		14'b10010100000011:	sigmoid = 21'b000000000000000000010;
		14'b10010100000100:	sigmoid = 21'b000000000000000000010;
		14'b10010100000101:	sigmoid = 21'b000000000000000000010;
		14'b10010100000110:	sigmoid = 21'b000000000000000000010;
		14'b10010100000111:	sigmoid = 21'b000000000000000000010;
		14'b10010100001000:	sigmoid = 21'b000000000000000000010;
		14'b10010100001001:	sigmoid = 21'b000000000000000000010;
		14'b10010100001010:	sigmoid = 21'b000000000000000000010;
		14'b10010100001011:	sigmoid = 21'b000000000000000000010;
		14'b10010100001100:	sigmoid = 21'b000000000000000000010;
		14'b10010100001101:	sigmoid = 21'b000000000000000000010;
		14'b10010100001110:	sigmoid = 21'b000000000000000000010;
		14'b10010100001111:	sigmoid = 21'b000000000000000000010;
		14'b10010100010000:	sigmoid = 21'b000000000000000000010;
		14'b10010100010001:	sigmoid = 21'b000000000000000000010;
		14'b10010100010010:	sigmoid = 21'b000000000000000000010;
		14'b10010100010011:	sigmoid = 21'b000000000000000000010;
		14'b10010100010100:	sigmoid = 21'b000000000000000000010;
		14'b10010100010101:	sigmoid = 21'b000000000000000000010;
		14'b10010100010110:	sigmoid = 21'b000000000000000000011;
		14'b10010100010111:	sigmoid = 21'b000000000000000000011;
		14'b10010100011000:	sigmoid = 21'b000000000000000000011;
		14'b10010100011001:	sigmoid = 21'b000000000000000000011;
		14'b10010100011010:	sigmoid = 21'b000000000000000000011;
		14'b10010100011011:	sigmoid = 21'b000000000000000000011;
		14'b10010100011100:	sigmoid = 21'b000000000000000000011;
		14'b10010100011101:	sigmoid = 21'b000000000000000000011;
		14'b10010100011110:	sigmoid = 21'b000000000000000000011;
		14'b10010100011111:	sigmoid = 21'b000000000000000000011;
		14'b10010100100000:	sigmoid = 21'b000000000000000000011;
		14'b10010100100001:	sigmoid = 21'b000000000000000000011;
		14'b10010100100010:	sigmoid = 21'b000000000000000000011;
		14'b10010100100011:	sigmoid = 21'b000000000000000000011;
		14'b10010100100100:	sigmoid = 21'b000000000000000000011;
		14'b10010100100101:	sigmoid = 21'b000000000000000000011;
		14'b10010100100110:	sigmoid = 21'b000000000000000000011;
		14'b10010100100111:	sigmoid = 21'b000000000000000000011;
		14'b10010100101000:	sigmoid = 21'b000000000000000000011;
		14'b10010100101001:	sigmoid = 21'b000000000000000000011;
		14'b10010100101010:	sigmoid = 21'b000000000000000000011;
		14'b10010100101011:	sigmoid = 21'b000000000000000000011;
		14'b10010100101100:	sigmoid = 21'b000000000000000000011;
		14'b10010100101101:	sigmoid = 21'b000000000000000000011;
		14'b10010100101110:	sigmoid = 21'b000000000000000000011;
		14'b10010100101111:	sigmoid = 21'b000000000000000000011;
		14'b10010100110000:	sigmoid = 21'b000000000000000000011;
		14'b10010100110001:	sigmoid = 21'b000000000000000000011;
		14'b10010100110010:	sigmoid = 21'b000000000000000000011;
		14'b10010100110011:	sigmoid = 21'b000000000000000000011;
		14'b10010100110100:	sigmoid = 21'b000000000000000000011;
		14'b10010100110101:	sigmoid = 21'b000000000000000000011;
		14'b10010100110110:	sigmoid = 21'b000000000000000000011;
		14'b10010100110111:	sigmoid = 21'b000000000000000000011;
		14'b10010100111000:	sigmoid = 21'b000000000000000000011;
		14'b10010100111001:	sigmoid = 21'b000000000000000000011;
		14'b10010100111010:	sigmoid = 21'b000000000000000000011;
		14'b10010100111011:	sigmoid = 21'b000000000000000000011;
		14'b10010100111100:	sigmoid = 21'b000000000000000000011;
		14'b10010100111101:	sigmoid = 21'b000000000000000000011;
		14'b10010100111110:	sigmoid = 21'b000000000000000000011;
		14'b10010100111111:	sigmoid = 21'b000000000000000000011;
		14'b10010101000000:	sigmoid = 21'b000000000000000000011;
		14'b10010101000001:	sigmoid = 21'b000000000000000000011;
		14'b10010101000010:	sigmoid = 21'b000000000000000000011;
		14'b10010101000011:	sigmoid = 21'b000000000000000000011;
		14'b10010101000100:	sigmoid = 21'b000000000000000000011;
		14'b10010101000101:	sigmoid = 21'b000000000000000000011;
		14'b10010101000110:	sigmoid = 21'b000000000000000000011;
		14'b10010101000111:	sigmoid = 21'b000000000000000000011;
		14'b10010101001000:	sigmoid = 21'b000000000000000000011;
		14'b10010101001001:	sigmoid = 21'b000000000000000000011;
		14'b10010101001010:	sigmoid = 21'b000000000000000000011;
		14'b10010101001011:	sigmoid = 21'b000000000000000000011;
		14'b10010101001100:	sigmoid = 21'b000000000000000000011;
		14'b10010101001101:	sigmoid = 21'b000000000000000000011;
		14'b10010101001110:	sigmoid = 21'b000000000000000000011;
		14'b10010101001111:	sigmoid = 21'b000000000000000000011;
		14'b10010101010000:	sigmoid = 21'b000000000000000000011;
		14'b10010101010001:	sigmoid = 21'b000000000000000000011;
		14'b10010101010010:	sigmoid = 21'b000000000000000000011;
		14'b10010101010011:	sigmoid = 21'b000000000000000000011;
		14'b10010101010100:	sigmoid = 21'b000000000000000000011;
		14'b10010101010101:	sigmoid = 21'b000000000000000000011;
		14'b10010101010110:	sigmoid = 21'b000000000000000000011;
		14'b10010101010111:	sigmoid = 21'b000000000000000000011;
		14'b10010101011000:	sigmoid = 21'b000000000000000000011;
		14'b10010101011001:	sigmoid = 21'b000000000000000000011;
		14'b10010101011010:	sigmoid = 21'b000000000000000000011;
		14'b10010101011011:	sigmoid = 21'b000000000000000000011;
		14'b10010101011100:	sigmoid = 21'b000000000000000000011;
		14'b10010101011101:	sigmoid = 21'b000000000000000000011;
		14'b10010101011110:	sigmoid = 21'b000000000000000000011;
		14'b10010101011111:	sigmoid = 21'b000000000000000000011;
		14'b10010101100000:	sigmoid = 21'b000000000000000000011;
		14'b10010101100001:	sigmoid = 21'b000000000000000000011;
		14'b10010101100010:	sigmoid = 21'b000000000000000000011;
		14'b10010101100011:	sigmoid = 21'b000000000000000000011;
		14'b10010101100100:	sigmoid = 21'b000000000000000000011;
		14'b10010101100101:	sigmoid = 21'b000000000000000000011;
		14'b10010101100110:	sigmoid = 21'b000000000000000000011;
		14'b10010101100111:	sigmoid = 21'b000000000000000000011;
		14'b10010101101000:	sigmoid = 21'b000000000000000000011;
		14'b10010101101001:	sigmoid = 21'b000000000000000000011;
		14'b10010101101010:	sigmoid = 21'b000000000000000000011;
		14'b10010101101011:	sigmoid = 21'b000000000000000000011;
		14'b10010101101100:	sigmoid = 21'b000000000000000000011;
		14'b10010101101101:	sigmoid = 21'b000000000000000000011;
		14'b10010101101110:	sigmoid = 21'b000000000000000000011;
		14'b10010101101111:	sigmoid = 21'b000000000000000000011;
		14'b10010101110000:	sigmoid = 21'b000000000000000000011;
		14'b10010101110001:	sigmoid = 21'b000000000000000000011;
		14'b10010101110010:	sigmoid = 21'b000000000000000000011;
		14'b10010101110011:	sigmoid = 21'b000000000000000000011;
		14'b10010101110100:	sigmoid = 21'b000000000000000000011;
		14'b10010101110101:	sigmoid = 21'b000000000000000000011;
		14'b10010101110110:	sigmoid = 21'b000000000000000000011;
		14'b10010101110111:	sigmoid = 21'b000000000000000000011;
		14'b10010101111000:	sigmoid = 21'b000000000000000000011;
		14'b10010101111001:	sigmoid = 21'b000000000000000000011;
		14'b10010101111010:	sigmoid = 21'b000000000000000000011;
		14'b10010101111011:	sigmoid = 21'b000000000000000000011;
		14'b10010101111100:	sigmoid = 21'b000000000000000000011;
		14'b10010101111101:	sigmoid = 21'b000000000000000000011;
		14'b10010101111110:	sigmoid = 21'b000000000000000000011;
		14'b10010101111111:	sigmoid = 21'b000000000000000000011;
		14'b10010110000000:	sigmoid = 21'b000000000000000000011;
		14'b10010110000001:	sigmoid = 21'b000000000000000000011;
		14'b10010110000010:	sigmoid = 21'b000000000000000000011;
		14'b10010110000011:	sigmoid = 21'b000000000000000000011;
		14'b10010110000100:	sigmoid = 21'b000000000000000000011;
		14'b10010110000101:	sigmoid = 21'b000000000000000000011;
		14'b10010110000110:	sigmoid = 21'b000000000000000000011;
		14'b10010110000111:	sigmoid = 21'b000000000000000000011;
		14'b10010110001000:	sigmoid = 21'b000000000000000000011;
		14'b10010110001001:	sigmoid = 21'b000000000000000000011;
		14'b10010110001010:	sigmoid = 21'b000000000000000000011;
		14'b10010110001011:	sigmoid = 21'b000000000000000000011;
		14'b10010110001100:	sigmoid = 21'b000000000000000000011;
		14'b10010110001101:	sigmoid = 21'b000000000000000000011;
		14'b10010110001110:	sigmoid = 21'b000000000000000000011;
		14'b10010110001111:	sigmoid = 21'b000000000000000000011;
		14'b10010110010000:	sigmoid = 21'b000000000000000000011;
		14'b10010110010001:	sigmoid = 21'b000000000000000000011;
		14'b10010110010010:	sigmoid = 21'b000000000000000000011;
		14'b10010110010011:	sigmoid = 21'b000000000000000000011;
		14'b10010110010100:	sigmoid = 21'b000000000000000000011;
		14'b10010110010101:	sigmoid = 21'b000000000000000000011;
		14'b10010110010110:	sigmoid = 21'b000000000000000000011;
		14'b10010110010111:	sigmoid = 21'b000000000000000000011;
		14'b10010110011000:	sigmoid = 21'b000000000000000000011;
		14'b10010110011001:	sigmoid = 21'b000000000000000000011;
		14'b10010110011010:	sigmoid = 21'b000000000000000000011;
		14'b10010110011011:	sigmoid = 21'b000000000000000000011;
		14'b10010110011100:	sigmoid = 21'b000000000000000000011;
		14'b10010110011101:	sigmoid = 21'b000000000000000000011;
		14'b10010110011110:	sigmoid = 21'b000000000000000000011;
		14'b10010110011111:	sigmoid = 21'b000000000000000000011;
		14'b10010110100000:	sigmoid = 21'b000000000000000000011;
		14'b10010110100001:	sigmoid = 21'b000000000000000000011;
		14'b10010110100010:	sigmoid = 21'b000000000000000000011;
		14'b10010110100011:	sigmoid = 21'b000000000000000000011;
		14'b10010110100100:	sigmoid = 21'b000000000000000000011;
		14'b10010110100101:	sigmoid = 21'b000000000000000000011;
		14'b10010110100110:	sigmoid = 21'b000000000000000000011;
		14'b10010110100111:	sigmoid = 21'b000000000000000000011;
		14'b10010110101000:	sigmoid = 21'b000000000000000000011;
		14'b10010110101001:	sigmoid = 21'b000000000000000000011;
		14'b10010110101010:	sigmoid = 21'b000000000000000000100;
		14'b10010110101011:	sigmoid = 21'b000000000000000000100;
		14'b10010110101100:	sigmoid = 21'b000000000000000000100;
		14'b10010110101101:	sigmoid = 21'b000000000000000000100;
		14'b10010110101110:	sigmoid = 21'b000000000000000000100;
		14'b10010110101111:	sigmoid = 21'b000000000000000000100;
		14'b10010110110000:	sigmoid = 21'b000000000000000000100;
		14'b10010110110001:	sigmoid = 21'b000000000000000000100;
		14'b10010110110010:	sigmoid = 21'b000000000000000000100;
		14'b10010110110011:	sigmoid = 21'b000000000000000000100;
		14'b10010110110100:	sigmoid = 21'b000000000000000000100;
		14'b10010110110101:	sigmoid = 21'b000000000000000000100;
		14'b10010110110110:	sigmoid = 21'b000000000000000000100;
		14'b10010110110111:	sigmoid = 21'b000000000000000000100;
		14'b10010110111000:	sigmoid = 21'b000000000000000000100;
		14'b10010110111001:	sigmoid = 21'b000000000000000000100;
		14'b10010110111010:	sigmoid = 21'b000000000000000000100;
		14'b10010110111011:	sigmoid = 21'b000000000000000000100;
		14'b10010110111100:	sigmoid = 21'b000000000000000000100;
		14'b10010110111101:	sigmoid = 21'b000000000000000000100;
		14'b10010110111110:	sigmoid = 21'b000000000000000000100;
		14'b10010110111111:	sigmoid = 21'b000000000000000000100;
		14'b10010111000000:	sigmoid = 21'b000000000000000000100;
		14'b10010111000001:	sigmoid = 21'b000000000000000000100;
		14'b10010111000010:	sigmoid = 21'b000000000000000000100;
		14'b10010111000011:	sigmoid = 21'b000000000000000000100;
		14'b10010111000100:	sigmoid = 21'b000000000000000000100;
		14'b10010111000101:	sigmoid = 21'b000000000000000000100;
		14'b10010111000110:	sigmoid = 21'b000000000000000000100;
		14'b10010111000111:	sigmoid = 21'b000000000000000000100;
		14'b10010111001000:	sigmoid = 21'b000000000000000000100;
		14'b10010111001001:	sigmoid = 21'b000000000000000000100;
		14'b10010111001010:	sigmoid = 21'b000000000000000000100;
		14'b10010111001011:	sigmoid = 21'b000000000000000000100;
		14'b10010111001100:	sigmoid = 21'b000000000000000000100;
		14'b10010111001101:	sigmoid = 21'b000000000000000000100;
		14'b10010111001110:	sigmoid = 21'b000000000000000000100;
		14'b10010111001111:	sigmoid = 21'b000000000000000000100;
		14'b10010111010000:	sigmoid = 21'b000000000000000000100;
		14'b10010111010001:	sigmoid = 21'b000000000000000000100;
		14'b10010111010010:	sigmoid = 21'b000000000000000000100;
		14'b10010111010011:	sigmoid = 21'b000000000000000000100;
		14'b10010111010100:	sigmoid = 21'b000000000000000000100;
		14'b10010111010101:	sigmoid = 21'b000000000000000000100;
		14'b10010111010110:	sigmoid = 21'b000000000000000000100;
		14'b10010111010111:	sigmoid = 21'b000000000000000000100;
		14'b10010111011000:	sigmoid = 21'b000000000000000000100;
		14'b10010111011001:	sigmoid = 21'b000000000000000000100;
		14'b10010111011010:	sigmoid = 21'b000000000000000000100;
		14'b10010111011011:	sigmoid = 21'b000000000000000000100;
		14'b10010111011100:	sigmoid = 21'b000000000000000000100;
		14'b10010111011101:	sigmoid = 21'b000000000000000000100;
		14'b10010111011110:	sigmoid = 21'b000000000000000000100;
		14'b10010111011111:	sigmoid = 21'b000000000000000000100;
		14'b10010111100000:	sigmoid = 21'b000000000000000000100;
		14'b10010111100001:	sigmoid = 21'b000000000000000000100;
		14'b10010111100010:	sigmoid = 21'b000000000000000000100;
		14'b10010111100011:	sigmoid = 21'b000000000000000000100;
		14'b10010111100100:	sigmoid = 21'b000000000000000000100;
		14'b10010111100101:	sigmoid = 21'b000000000000000000100;
		14'b10010111100110:	sigmoid = 21'b000000000000000000100;
		14'b10010111100111:	sigmoid = 21'b000000000000000000100;
		14'b10010111101000:	sigmoid = 21'b000000000000000000100;
		14'b10010111101001:	sigmoid = 21'b000000000000000000100;
		14'b10010111101010:	sigmoid = 21'b000000000000000000100;
		14'b10010111101011:	sigmoid = 21'b000000000000000000100;
		14'b10010111101100:	sigmoid = 21'b000000000000000000100;
		14'b10010111101101:	sigmoid = 21'b000000000000000000100;
		14'b10010111101110:	sigmoid = 21'b000000000000000000100;
		14'b10010111101111:	sigmoid = 21'b000000000000000000100;
		14'b10010111110000:	sigmoid = 21'b000000000000000000100;
		14'b10010111110001:	sigmoid = 21'b000000000000000000100;
		14'b10010111110010:	sigmoid = 21'b000000000000000000100;
		14'b10010111110011:	sigmoid = 21'b000000000000000000100;
		14'b10010111110100:	sigmoid = 21'b000000000000000000100;
		14'b10010111110101:	sigmoid = 21'b000000000000000000100;
		14'b10010111110110:	sigmoid = 21'b000000000000000000100;
		14'b10010111110111:	sigmoid = 21'b000000000000000000100;
		14'b10010111111000:	sigmoid = 21'b000000000000000000100;
		14'b10010111111001:	sigmoid = 21'b000000000000000000100;
		14'b10010111111010:	sigmoid = 21'b000000000000000000100;
		14'b10010111111011:	sigmoid = 21'b000000000000000000100;
		14'b10010111111100:	sigmoid = 21'b000000000000000000100;
		14'b10010111111101:	sigmoid = 21'b000000000000000000100;
		14'b10010111111110:	sigmoid = 21'b000000000000000000100;
		14'b10010111111111:	sigmoid = 21'b000000000000000000100;
		14'b10011000000000:	sigmoid = 21'b000000000000000000100;
		14'b10011000000001:	sigmoid = 21'b000000000000000000100;
		14'b10011000000010:	sigmoid = 21'b000000000000000000100;
		14'b10011000000011:	sigmoid = 21'b000000000000000000100;
		14'b10011000000100:	sigmoid = 21'b000000000000000000100;
		14'b10011000000101:	sigmoid = 21'b000000000000000000100;
		14'b10011000000110:	sigmoid = 21'b000000000000000000100;
		14'b10011000000111:	sigmoid = 21'b000000000000000000100;
		14'b10011000001000:	sigmoid = 21'b000000000000000000100;
		14'b10011000001001:	sigmoid = 21'b000000000000000000100;
		14'b10011000001010:	sigmoid = 21'b000000000000000000100;
		14'b10011000001011:	sigmoid = 21'b000000000000000000100;
		14'b10011000001100:	sigmoid = 21'b000000000000000000100;
		14'b10011000001101:	sigmoid = 21'b000000000000000000100;
		14'b10011000001110:	sigmoid = 21'b000000000000000000100;
		14'b10011000001111:	sigmoid = 21'b000000000000000000100;
		14'b10011000010000:	sigmoid = 21'b000000000000000000100;
		14'b10011000010001:	sigmoid = 21'b000000000000000000100;
		14'b10011000010010:	sigmoid = 21'b000000000000000000100;
		14'b10011000010011:	sigmoid = 21'b000000000000000000100;
		14'b10011000010100:	sigmoid = 21'b000000000000000000100;
		14'b10011000010101:	sigmoid = 21'b000000000000000000100;
		14'b10011000010110:	sigmoid = 21'b000000000000000000100;
		14'b10011000010111:	sigmoid = 21'b000000000000000000100;
		14'b10011000011000:	sigmoid = 21'b000000000000000000100;
		14'b10011000011001:	sigmoid = 21'b000000000000000000100;
		14'b10011000011010:	sigmoid = 21'b000000000000000000100;
		14'b10011000011011:	sigmoid = 21'b000000000000000000100;
		14'b10011000011100:	sigmoid = 21'b000000000000000000101;
		14'b10011000011101:	sigmoid = 21'b000000000000000000101;
		14'b10011000011110:	sigmoid = 21'b000000000000000000101;
		14'b10011000011111:	sigmoid = 21'b000000000000000000101;
		14'b10011000100000:	sigmoid = 21'b000000000000000000101;
		14'b10011000100001:	sigmoid = 21'b000000000000000000101;
		14'b10011000100010:	sigmoid = 21'b000000000000000000101;
		14'b10011000100011:	sigmoid = 21'b000000000000000000101;
		14'b10011000100100:	sigmoid = 21'b000000000000000000101;
		14'b10011000100101:	sigmoid = 21'b000000000000000000101;
		14'b10011000100110:	sigmoid = 21'b000000000000000000101;
		14'b10011000100111:	sigmoid = 21'b000000000000000000101;
		14'b10011000101000:	sigmoid = 21'b000000000000000000101;
		14'b10011000101001:	sigmoid = 21'b000000000000000000101;
		14'b10011000101010:	sigmoid = 21'b000000000000000000101;
		14'b10011000101011:	sigmoid = 21'b000000000000000000101;
		14'b10011000101100:	sigmoid = 21'b000000000000000000101;
		14'b10011000101101:	sigmoid = 21'b000000000000000000101;
		14'b10011000101110:	sigmoid = 21'b000000000000000000101;
		14'b10011000101111:	sigmoid = 21'b000000000000000000101;
		14'b10011000110000:	sigmoid = 21'b000000000000000000101;
		14'b10011000110001:	sigmoid = 21'b000000000000000000101;
		14'b10011000110010:	sigmoid = 21'b000000000000000000101;
		14'b10011000110011:	sigmoid = 21'b000000000000000000101;
		14'b10011000110100:	sigmoid = 21'b000000000000000000101;
		14'b10011000110101:	sigmoid = 21'b000000000000000000101;
		14'b10011000110110:	sigmoid = 21'b000000000000000000101;
		14'b10011000110111:	sigmoid = 21'b000000000000000000101;
		14'b10011000111000:	sigmoid = 21'b000000000000000000101;
		14'b10011000111001:	sigmoid = 21'b000000000000000000101;
		14'b10011000111010:	sigmoid = 21'b000000000000000000101;
		14'b10011000111011:	sigmoid = 21'b000000000000000000101;
		14'b10011000111100:	sigmoid = 21'b000000000000000000101;
		14'b10011000111101:	sigmoid = 21'b000000000000000000101;
		14'b10011000111110:	sigmoid = 21'b000000000000000000101;
		14'b10011000111111:	sigmoid = 21'b000000000000000000101;
		14'b10011001000000:	sigmoid = 21'b000000000000000000101;
		14'b10011001000001:	sigmoid = 21'b000000000000000000101;
		14'b10011001000010:	sigmoid = 21'b000000000000000000101;
		14'b10011001000011:	sigmoid = 21'b000000000000000000101;
		14'b10011001000100:	sigmoid = 21'b000000000000000000101;
		14'b10011001000101:	sigmoid = 21'b000000000000000000101;
		14'b10011001000110:	sigmoid = 21'b000000000000000000101;
		14'b10011001000111:	sigmoid = 21'b000000000000000000101;
		14'b10011001001000:	sigmoid = 21'b000000000000000000101;
		14'b10011001001001:	sigmoid = 21'b000000000000000000101;
		14'b10011001001010:	sigmoid = 21'b000000000000000000101;
		14'b10011001001011:	sigmoid = 21'b000000000000000000101;
		14'b10011001001100:	sigmoid = 21'b000000000000000000101;
		14'b10011001001101:	sigmoid = 21'b000000000000000000101;
		14'b10011001001110:	sigmoid = 21'b000000000000000000101;
		14'b10011001001111:	sigmoid = 21'b000000000000000000101;
		14'b10011001010000:	sigmoid = 21'b000000000000000000101;
		14'b10011001010001:	sigmoid = 21'b000000000000000000101;
		14'b10011001010010:	sigmoid = 21'b000000000000000000101;
		14'b10011001010011:	sigmoid = 21'b000000000000000000101;
		14'b10011001010100:	sigmoid = 21'b000000000000000000101;
		14'b10011001010101:	sigmoid = 21'b000000000000000000101;
		14'b10011001010110:	sigmoid = 21'b000000000000000000101;
		14'b10011001010111:	sigmoid = 21'b000000000000000000101;
		14'b10011001011000:	sigmoid = 21'b000000000000000000101;
		14'b10011001011001:	sigmoid = 21'b000000000000000000101;
		14'b10011001011010:	sigmoid = 21'b000000000000000000101;
		14'b10011001011011:	sigmoid = 21'b000000000000000000101;
		14'b10011001011100:	sigmoid = 21'b000000000000000000101;
		14'b10011001011101:	sigmoid = 21'b000000000000000000101;
		14'b10011001011110:	sigmoid = 21'b000000000000000000101;
		14'b10011001011111:	sigmoid = 21'b000000000000000000101;
		14'b10011001100000:	sigmoid = 21'b000000000000000000101;
		14'b10011001100001:	sigmoid = 21'b000000000000000000101;
		14'b10011001100010:	sigmoid = 21'b000000000000000000101;
		14'b10011001100011:	sigmoid = 21'b000000000000000000101;
		14'b10011001100100:	sigmoid = 21'b000000000000000000101;
		14'b10011001100101:	sigmoid = 21'b000000000000000000101;
		14'b10011001100110:	sigmoid = 21'b000000000000000000101;
		14'b10011001100111:	sigmoid = 21'b000000000000000000101;
		14'b10011001101000:	sigmoid = 21'b000000000000000000101;
		14'b10011001101001:	sigmoid = 21'b000000000000000000101;
		14'b10011001101010:	sigmoid = 21'b000000000000000000101;
		14'b10011001101011:	sigmoid = 21'b000000000000000000101;
		14'b10011001101100:	sigmoid = 21'b000000000000000000101;
		14'b10011001101101:	sigmoid = 21'b000000000000000000101;
		14'b10011001101110:	sigmoid = 21'b000000000000000000101;
		14'b10011001101111:	sigmoid = 21'b000000000000000000101;
		14'b10011001110000:	sigmoid = 21'b000000000000000000101;
		14'b10011001110001:	sigmoid = 21'b000000000000000000101;
		14'b10011001110010:	sigmoid = 21'b000000000000000000101;
		14'b10011001110011:	sigmoid = 21'b000000000000000000101;
		14'b10011001110100:	sigmoid = 21'b000000000000000000101;
		14'b10011001110101:	sigmoid = 21'b000000000000000000101;
		14'b10011001110110:	sigmoid = 21'b000000000000000000101;
		14'b10011001110111:	sigmoid = 21'b000000000000000000101;
		14'b10011001111000:	sigmoid = 21'b000000000000000000101;
		14'b10011001111001:	sigmoid = 21'b000000000000000000110;
		14'b10011001111010:	sigmoid = 21'b000000000000000000110;
		14'b10011001111011:	sigmoid = 21'b000000000000000000110;
		14'b10011001111100:	sigmoid = 21'b000000000000000000110;
		14'b10011001111101:	sigmoid = 21'b000000000000000000110;
		14'b10011001111110:	sigmoid = 21'b000000000000000000110;
		14'b10011001111111:	sigmoid = 21'b000000000000000000110;
		14'b10011010000000:	sigmoid = 21'b000000000000000000110;
		14'b10011010000001:	sigmoid = 21'b000000000000000000110;
		14'b10011010000010:	sigmoid = 21'b000000000000000000110;
		14'b10011010000011:	sigmoid = 21'b000000000000000000110;
		14'b10011010000100:	sigmoid = 21'b000000000000000000110;
		14'b10011010000101:	sigmoid = 21'b000000000000000000110;
		14'b10011010000110:	sigmoid = 21'b000000000000000000110;
		14'b10011010000111:	sigmoid = 21'b000000000000000000110;
		14'b10011010001000:	sigmoid = 21'b000000000000000000110;
		14'b10011010001001:	sigmoid = 21'b000000000000000000110;
		14'b10011010001010:	sigmoid = 21'b000000000000000000110;
		14'b10011010001011:	sigmoid = 21'b000000000000000000110;
		14'b10011010001100:	sigmoid = 21'b000000000000000000110;
		14'b10011010001101:	sigmoid = 21'b000000000000000000110;
		14'b10011010001110:	sigmoid = 21'b000000000000000000110;
		14'b10011010001111:	sigmoid = 21'b000000000000000000110;
		14'b10011010010000:	sigmoid = 21'b000000000000000000110;
		14'b10011010010001:	sigmoid = 21'b000000000000000000110;
		14'b10011010010010:	sigmoid = 21'b000000000000000000110;
		14'b10011010010011:	sigmoid = 21'b000000000000000000110;
		14'b10011010010100:	sigmoid = 21'b000000000000000000110;
		14'b10011010010101:	sigmoid = 21'b000000000000000000110;
		14'b10011010010110:	sigmoid = 21'b000000000000000000110;
		14'b10011010010111:	sigmoid = 21'b000000000000000000110;
		14'b10011010011000:	sigmoid = 21'b000000000000000000110;
		14'b10011010011001:	sigmoid = 21'b000000000000000000110;
		14'b10011010011010:	sigmoid = 21'b000000000000000000110;
		14'b10011010011011:	sigmoid = 21'b000000000000000000110;
		14'b10011010011100:	sigmoid = 21'b000000000000000000110;
		14'b10011010011101:	sigmoid = 21'b000000000000000000110;
		14'b10011010011110:	sigmoid = 21'b000000000000000000110;
		14'b10011010011111:	sigmoid = 21'b000000000000000000110;
		14'b10011010100000:	sigmoid = 21'b000000000000000000110;
		14'b10011010100001:	sigmoid = 21'b000000000000000000110;
		14'b10011010100010:	sigmoid = 21'b000000000000000000110;
		14'b10011010100011:	sigmoid = 21'b000000000000000000110;
		14'b10011010100100:	sigmoid = 21'b000000000000000000110;
		14'b10011010100101:	sigmoid = 21'b000000000000000000110;
		14'b10011010100110:	sigmoid = 21'b000000000000000000110;
		14'b10011010100111:	sigmoid = 21'b000000000000000000110;
		14'b10011010101000:	sigmoid = 21'b000000000000000000110;
		14'b10011010101001:	sigmoid = 21'b000000000000000000110;
		14'b10011010101010:	sigmoid = 21'b000000000000000000110;
		14'b10011010101011:	sigmoid = 21'b000000000000000000110;
		14'b10011010101100:	sigmoid = 21'b000000000000000000110;
		14'b10011010101101:	sigmoid = 21'b000000000000000000110;
		14'b10011010101110:	sigmoid = 21'b000000000000000000110;
		14'b10011010101111:	sigmoid = 21'b000000000000000000110;
		14'b10011010110000:	sigmoid = 21'b000000000000000000110;
		14'b10011010110001:	sigmoid = 21'b000000000000000000110;
		14'b10011010110010:	sigmoid = 21'b000000000000000000110;
		14'b10011010110011:	sigmoid = 21'b000000000000000000110;
		14'b10011010110100:	sigmoid = 21'b000000000000000000110;
		14'b10011010110101:	sigmoid = 21'b000000000000000000110;
		14'b10011010110110:	sigmoid = 21'b000000000000000000110;
		14'b10011010110111:	sigmoid = 21'b000000000000000000110;
		14'b10011010111000:	sigmoid = 21'b000000000000000000110;
		14'b10011010111001:	sigmoid = 21'b000000000000000000110;
		14'b10011010111010:	sigmoid = 21'b000000000000000000110;
		14'b10011010111011:	sigmoid = 21'b000000000000000000110;
		14'b10011010111100:	sigmoid = 21'b000000000000000000110;
		14'b10011010111101:	sigmoid = 21'b000000000000000000110;
		14'b10011010111110:	sigmoid = 21'b000000000000000000110;
		14'b10011010111111:	sigmoid = 21'b000000000000000000110;
		14'b10011011000000:	sigmoid = 21'b000000000000000000110;
		14'b10011011000001:	sigmoid = 21'b000000000000000000110;
		14'b10011011000010:	sigmoid = 21'b000000000000000000110;
		14'b10011011000011:	sigmoid = 21'b000000000000000000110;
		14'b10011011000100:	sigmoid = 21'b000000000000000000110;
		14'b10011011000101:	sigmoid = 21'b000000000000000000110;
		14'b10011011000110:	sigmoid = 21'b000000000000000000110;
		14'b10011011000111:	sigmoid = 21'b000000000000000000110;
		14'b10011011001000:	sigmoid = 21'b000000000000000000111;
		14'b10011011001001:	sigmoid = 21'b000000000000000000111;
		14'b10011011001010:	sigmoid = 21'b000000000000000000111;
		14'b10011011001011:	sigmoid = 21'b000000000000000000111;
		14'b10011011001100:	sigmoid = 21'b000000000000000000111;
		14'b10011011001101:	sigmoid = 21'b000000000000000000111;
		14'b10011011001110:	sigmoid = 21'b000000000000000000111;
		14'b10011011001111:	sigmoid = 21'b000000000000000000111;
		14'b10011011010000:	sigmoid = 21'b000000000000000000111;
		14'b10011011010001:	sigmoid = 21'b000000000000000000111;
		14'b10011011010010:	sigmoid = 21'b000000000000000000111;
		14'b10011011010011:	sigmoid = 21'b000000000000000000111;
		14'b10011011010100:	sigmoid = 21'b000000000000000000111;
		14'b10011011010101:	sigmoid = 21'b000000000000000000111;
		14'b10011011010110:	sigmoid = 21'b000000000000000000111;
		14'b10011011010111:	sigmoid = 21'b000000000000000000111;
		14'b10011011011000:	sigmoid = 21'b000000000000000000111;
		14'b10011011011001:	sigmoid = 21'b000000000000000000111;
		14'b10011011011010:	sigmoid = 21'b000000000000000000111;
		14'b10011011011011:	sigmoid = 21'b000000000000000000111;
		14'b10011011011100:	sigmoid = 21'b000000000000000000111;
		14'b10011011011101:	sigmoid = 21'b000000000000000000111;
		14'b10011011011110:	sigmoid = 21'b000000000000000000111;
		14'b10011011011111:	sigmoid = 21'b000000000000000000111;
		14'b10011011100000:	sigmoid = 21'b000000000000000000111;
		14'b10011011100001:	sigmoid = 21'b000000000000000000111;
		14'b10011011100010:	sigmoid = 21'b000000000000000000111;
		14'b10011011100011:	sigmoid = 21'b000000000000000000111;
		14'b10011011100100:	sigmoid = 21'b000000000000000000111;
		14'b10011011100101:	sigmoid = 21'b000000000000000000111;
		14'b10011011100110:	sigmoid = 21'b000000000000000000111;
		14'b10011011100111:	sigmoid = 21'b000000000000000000111;
		14'b10011011101000:	sigmoid = 21'b000000000000000000111;
		14'b10011011101001:	sigmoid = 21'b000000000000000000111;
		14'b10011011101010:	sigmoid = 21'b000000000000000000111;
		14'b10011011101011:	sigmoid = 21'b000000000000000000111;
		14'b10011011101100:	sigmoid = 21'b000000000000000000111;
		14'b10011011101101:	sigmoid = 21'b000000000000000000111;
		14'b10011011101110:	sigmoid = 21'b000000000000000000111;
		14'b10011011101111:	sigmoid = 21'b000000000000000000111;
		14'b10011011110000:	sigmoid = 21'b000000000000000000111;
		14'b10011011110001:	sigmoid = 21'b000000000000000000111;
		14'b10011011110010:	sigmoid = 21'b000000000000000000111;
		14'b10011011110011:	sigmoid = 21'b000000000000000000111;
		14'b10011011110100:	sigmoid = 21'b000000000000000000111;
		14'b10011011110101:	sigmoid = 21'b000000000000000000111;
		14'b10011011110110:	sigmoid = 21'b000000000000000000111;
		14'b10011011110111:	sigmoid = 21'b000000000000000000111;
		14'b10011011111000:	sigmoid = 21'b000000000000000000111;
		14'b10011011111001:	sigmoid = 21'b000000000000000000111;
		14'b10011011111010:	sigmoid = 21'b000000000000000000111;
		14'b10011011111011:	sigmoid = 21'b000000000000000000111;
		14'b10011011111100:	sigmoid = 21'b000000000000000000111;
		14'b10011011111101:	sigmoid = 21'b000000000000000000111;
		14'b10011011111110:	sigmoid = 21'b000000000000000000111;
		14'b10011011111111:	sigmoid = 21'b000000000000000000111;
		14'b10011100000000:	sigmoid = 21'b000000000000000000111;
		14'b10011100000001:	sigmoid = 21'b000000000000000000111;
		14'b10011100000010:	sigmoid = 21'b000000000000000000111;
		14'b10011100000011:	sigmoid = 21'b000000000000000000111;
		14'b10011100000100:	sigmoid = 21'b000000000000000000111;
		14'b10011100000101:	sigmoid = 21'b000000000000000000111;
		14'b10011100000110:	sigmoid = 21'b000000000000000000111;
		14'b10011100000111:	sigmoid = 21'b000000000000000000111;
		14'b10011100001000:	sigmoid = 21'b000000000000000000111;
		14'b10011100001001:	sigmoid = 21'b000000000000000000111;
		14'b10011100001010:	sigmoid = 21'b000000000000000000111;
		14'b10011100001011:	sigmoid = 21'b000000000000000000111;
		14'b10011100001100:	sigmoid = 21'b000000000000000001000;
		14'b10011100001101:	sigmoid = 21'b000000000000000001000;
		14'b10011100001110:	sigmoid = 21'b000000000000000001000;
		14'b10011100001111:	sigmoid = 21'b000000000000000001000;
		14'b10011100010000:	sigmoid = 21'b000000000000000001000;
		14'b10011100010001:	sigmoid = 21'b000000000000000001000;
		14'b10011100010010:	sigmoid = 21'b000000000000000001000;
		14'b10011100010011:	sigmoid = 21'b000000000000000001000;
		14'b10011100010100:	sigmoid = 21'b000000000000000001000;
		14'b10011100010101:	sigmoid = 21'b000000000000000001000;
		14'b10011100010110:	sigmoid = 21'b000000000000000001000;
		14'b10011100010111:	sigmoid = 21'b000000000000000001000;
		14'b10011100011000:	sigmoid = 21'b000000000000000001000;
		14'b10011100011001:	sigmoid = 21'b000000000000000001000;
		14'b10011100011010:	sigmoid = 21'b000000000000000001000;
		14'b10011100011011:	sigmoid = 21'b000000000000000001000;
		14'b10011100011100:	sigmoid = 21'b000000000000000001000;
		14'b10011100011101:	sigmoid = 21'b000000000000000001000;
		14'b10011100011110:	sigmoid = 21'b000000000000000001000;
		14'b10011100011111:	sigmoid = 21'b000000000000000001000;
		14'b10011100100000:	sigmoid = 21'b000000000000000001000;
		14'b10011100100001:	sigmoid = 21'b000000000000000001000;
		14'b10011100100010:	sigmoid = 21'b000000000000000001000;
		14'b10011100100011:	sigmoid = 21'b000000000000000001000;
		14'b10011100100100:	sigmoid = 21'b000000000000000001000;
		14'b10011100100101:	sigmoid = 21'b000000000000000001000;
		14'b10011100100110:	sigmoid = 21'b000000000000000001000;
		14'b10011100100111:	sigmoid = 21'b000000000000000001000;
		14'b10011100101000:	sigmoid = 21'b000000000000000001000;
		14'b10011100101001:	sigmoid = 21'b000000000000000001000;
		14'b10011100101010:	sigmoid = 21'b000000000000000001000;
		14'b10011100101011:	sigmoid = 21'b000000000000000001000;
		14'b10011100101100:	sigmoid = 21'b000000000000000001000;
		14'b10011100101101:	sigmoid = 21'b000000000000000001000;
		14'b10011100101110:	sigmoid = 21'b000000000000000001000;
		14'b10011100101111:	sigmoid = 21'b000000000000000001000;
		14'b10011100110000:	sigmoid = 21'b000000000000000001000;
		14'b10011100110001:	sigmoid = 21'b000000000000000001000;
		14'b10011100110010:	sigmoid = 21'b000000000000000001000;
		14'b10011100110011:	sigmoid = 21'b000000000000000001000;
		14'b10011100110100:	sigmoid = 21'b000000000000000001000;
		14'b10011100110101:	sigmoid = 21'b000000000000000001000;
		14'b10011100110110:	sigmoid = 21'b000000000000000001000;
		14'b10011100110111:	sigmoid = 21'b000000000000000001000;
		14'b10011100111000:	sigmoid = 21'b000000000000000001000;
		14'b10011100111001:	sigmoid = 21'b000000000000000001000;
		14'b10011100111010:	sigmoid = 21'b000000000000000001000;
		14'b10011100111011:	sigmoid = 21'b000000000000000001000;
		14'b10011100111100:	sigmoid = 21'b000000000000000001000;
		14'b10011100111101:	sigmoid = 21'b000000000000000001000;
		14'b10011100111110:	sigmoid = 21'b000000000000000001000;
		14'b10011100111111:	sigmoid = 21'b000000000000000001000;
		14'b10011101000000:	sigmoid = 21'b000000000000000001000;
		14'b10011101000001:	sigmoid = 21'b000000000000000001000;
		14'b10011101000010:	sigmoid = 21'b000000000000000001000;
		14'b10011101000011:	sigmoid = 21'b000000000000000001000;
		14'b10011101000100:	sigmoid = 21'b000000000000000001000;
		14'b10011101000101:	sigmoid = 21'b000000000000000001000;
		14'b10011101000110:	sigmoid = 21'b000000000000000001000;
		14'b10011101000111:	sigmoid = 21'b000000000000000001000;
		14'b10011101001000:	sigmoid = 21'b000000000000000001000;
		14'b10011101001001:	sigmoid = 21'b000000000000000001001;
		14'b10011101001010:	sigmoid = 21'b000000000000000001001;
		14'b10011101001011:	sigmoid = 21'b000000000000000001001;
		14'b10011101001100:	sigmoid = 21'b000000000000000001001;
		14'b10011101001101:	sigmoid = 21'b000000000000000001001;
		14'b10011101001110:	sigmoid = 21'b000000000000000001001;
		14'b10011101001111:	sigmoid = 21'b000000000000000001001;
		14'b10011101010000:	sigmoid = 21'b000000000000000001001;
		14'b10011101010001:	sigmoid = 21'b000000000000000001001;
		14'b10011101010010:	sigmoid = 21'b000000000000000001001;
		14'b10011101010011:	sigmoid = 21'b000000000000000001001;
		14'b10011101010100:	sigmoid = 21'b000000000000000001001;
		14'b10011101010101:	sigmoid = 21'b000000000000000001001;
		14'b10011101010110:	sigmoid = 21'b000000000000000001001;
		14'b10011101010111:	sigmoid = 21'b000000000000000001001;
		14'b10011101011000:	sigmoid = 21'b000000000000000001001;
		14'b10011101011001:	sigmoid = 21'b000000000000000001001;
		14'b10011101011010:	sigmoid = 21'b000000000000000001001;
		14'b10011101011011:	sigmoid = 21'b000000000000000001001;
		14'b10011101011100:	sigmoid = 21'b000000000000000001001;
		14'b10011101011101:	sigmoid = 21'b000000000000000001001;
		14'b10011101011110:	sigmoid = 21'b000000000000000001001;
		14'b10011101011111:	sigmoid = 21'b000000000000000001001;
		14'b10011101100000:	sigmoid = 21'b000000000000000001001;
		14'b10011101100001:	sigmoid = 21'b000000000000000001001;
		14'b10011101100010:	sigmoid = 21'b000000000000000001001;
		14'b10011101100011:	sigmoid = 21'b000000000000000001001;
		14'b10011101100100:	sigmoid = 21'b000000000000000001001;
		14'b10011101100101:	sigmoid = 21'b000000000000000001001;
		14'b10011101100110:	sigmoid = 21'b000000000000000001001;
		14'b10011101100111:	sigmoid = 21'b000000000000000001001;
		14'b10011101101000:	sigmoid = 21'b000000000000000001001;
		14'b10011101101001:	sigmoid = 21'b000000000000000001001;
		14'b10011101101010:	sigmoid = 21'b000000000000000001001;
		14'b10011101101011:	sigmoid = 21'b000000000000000001001;
		14'b10011101101100:	sigmoid = 21'b000000000000000001001;
		14'b10011101101101:	sigmoid = 21'b000000000000000001001;
		14'b10011101101110:	sigmoid = 21'b000000000000000001001;
		14'b10011101101111:	sigmoid = 21'b000000000000000001001;
		14'b10011101110000:	sigmoid = 21'b000000000000000001001;
		14'b10011101110001:	sigmoid = 21'b000000000000000001001;
		14'b10011101110010:	sigmoid = 21'b000000000000000001001;
		14'b10011101110011:	sigmoid = 21'b000000000000000001001;
		14'b10011101110100:	sigmoid = 21'b000000000000000001001;
		14'b10011101110101:	sigmoid = 21'b000000000000000001001;
		14'b10011101110110:	sigmoid = 21'b000000000000000001001;
		14'b10011101110111:	sigmoid = 21'b000000000000000001001;
		14'b10011101111000:	sigmoid = 21'b000000000000000001001;
		14'b10011101111001:	sigmoid = 21'b000000000000000001001;
		14'b10011101111010:	sigmoid = 21'b000000000000000001001;
		14'b10011101111011:	sigmoid = 21'b000000000000000001001;
		14'b10011101111100:	sigmoid = 21'b000000000000000001001;
		14'b10011101111101:	sigmoid = 21'b000000000000000001001;
		14'b10011101111110:	sigmoid = 21'b000000000000000001001;
		14'b10011101111111:	sigmoid = 21'b000000000000000001010;
		14'b10011110000000:	sigmoid = 21'b000000000000000001010;
		14'b10011110000001:	sigmoid = 21'b000000000000000001010;
		14'b10011110000010:	sigmoid = 21'b000000000000000001010;
		14'b10011110000011:	sigmoid = 21'b000000000000000001010;
		14'b10011110000100:	sigmoid = 21'b000000000000000001010;
		14'b10011110000101:	sigmoid = 21'b000000000000000001010;
		14'b10011110000110:	sigmoid = 21'b000000000000000001010;
		14'b10011110000111:	sigmoid = 21'b000000000000000001010;
		14'b10011110001000:	sigmoid = 21'b000000000000000001010;
		14'b10011110001001:	sigmoid = 21'b000000000000000001010;
		14'b10011110001010:	sigmoid = 21'b000000000000000001010;
		14'b10011110001011:	sigmoid = 21'b000000000000000001010;
		14'b10011110001100:	sigmoid = 21'b000000000000000001010;
		14'b10011110001101:	sigmoid = 21'b000000000000000001010;
		14'b10011110001110:	sigmoid = 21'b000000000000000001010;
		14'b10011110001111:	sigmoid = 21'b000000000000000001010;
		14'b10011110010000:	sigmoid = 21'b000000000000000001010;
		14'b10011110010001:	sigmoid = 21'b000000000000000001010;
		14'b10011110010010:	sigmoid = 21'b000000000000000001010;
		14'b10011110010011:	sigmoid = 21'b000000000000000001010;
		14'b10011110010100:	sigmoid = 21'b000000000000000001010;
		14'b10011110010101:	sigmoid = 21'b000000000000000001010;
		14'b10011110010110:	sigmoid = 21'b000000000000000001010;
		14'b10011110010111:	sigmoid = 21'b000000000000000001010;
		14'b10011110011000:	sigmoid = 21'b000000000000000001010;
		14'b10011110011001:	sigmoid = 21'b000000000000000001010;
		14'b10011110011010:	sigmoid = 21'b000000000000000001010;
		14'b10011110011011:	sigmoid = 21'b000000000000000001010;
		14'b10011110011100:	sigmoid = 21'b000000000000000001010;
		14'b10011110011101:	sigmoid = 21'b000000000000000001010;
		14'b10011110011110:	sigmoid = 21'b000000000000000001010;
		14'b10011110011111:	sigmoid = 21'b000000000000000001010;
		14'b10011110100000:	sigmoid = 21'b000000000000000001010;
		14'b10011110100001:	sigmoid = 21'b000000000000000001010;
		14'b10011110100010:	sigmoid = 21'b000000000000000001010;
		14'b10011110100011:	sigmoid = 21'b000000000000000001010;
		14'b10011110100100:	sigmoid = 21'b000000000000000001010;
		14'b10011110100101:	sigmoid = 21'b000000000000000001010;
		14'b10011110100110:	sigmoid = 21'b000000000000000001010;
		14'b10011110100111:	sigmoid = 21'b000000000000000001010;
		14'b10011110101000:	sigmoid = 21'b000000000000000001010;
		14'b10011110101001:	sigmoid = 21'b000000000000000001010;
		14'b10011110101010:	sigmoid = 21'b000000000000000001010;
		14'b10011110101011:	sigmoid = 21'b000000000000000001010;
		14'b10011110101100:	sigmoid = 21'b000000000000000001010;
		14'b10011110101101:	sigmoid = 21'b000000000000000001010;
		14'b10011110101110:	sigmoid = 21'b000000000000000001010;
		14'b10011110101111:	sigmoid = 21'b000000000000000001010;
		14'b10011110110000:	sigmoid = 21'b000000000000000001011;
		14'b10011110110001:	sigmoid = 21'b000000000000000001011;
		14'b10011110110010:	sigmoid = 21'b000000000000000001011;
		14'b10011110110011:	sigmoid = 21'b000000000000000001011;
		14'b10011110110100:	sigmoid = 21'b000000000000000001011;
		14'b10011110110101:	sigmoid = 21'b000000000000000001011;
		14'b10011110110110:	sigmoid = 21'b000000000000000001011;
		14'b10011110110111:	sigmoid = 21'b000000000000000001011;
		14'b10011110111000:	sigmoid = 21'b000000000000000001011;
		14'b10011110111001:	sigmoid = 21'b000000000000000001011;
		14'b10011110111010:	sigmoid = 21'b000000000000000001011;
		14'b10011110111011:	sigmoid = 21'b000000000000000001011;
		14'b10011110111100:	sigmoid = 21'b000000000000000001011;
		14'b10011110111101:	sigmoid = 21'b000000000000000001011;
		14'b10011110111110:	sigmoid = 21'b000000000000000001011;
		14'b10011110111111:	sigmoid = 21'b000000000000000001011;
		14'b10011111000000:	sigmoid = 21'b000000000000000001011;
		14'b10011111000001:	sigmoid = 21'b000000000000000001011;
		14'b10011111000010:	sigmoid = 21'b000000000000000001011;
		14'b10011111000011:	sigmoid = 21'b000000000000000001011;
		14'b10011111000100:	sigmoid = 21'b000000000000000001011;
		14'b10011111000101:	sigmoid = 21'b000000000000000001011;
		14'b10011111000110:	sigmoid = 21'b000000000000000001011;
		14'b10011111000111:	sigmoid = 21'b000000000000000001011;
		14'b10011111001000:	sigmoid = 21'b000000000000000001011;
		14'b10011111001001:	sigmoid = 21'b000000000000000001011;
		14'b10011111001010:	sigmoid = 21'b000000000000000001011;
		14'b10011111001011:	sigmoid = 21'b000000000000000001011;
		14'b10011111001100:	sigmoid = 21'b000000000000000001011;
		14'b10011111001101:	sigmoid = 21'b000000000000000001011;
		14'b10011111001110:	sigmoid = 21'b000000000000000001011;
		14'b10011111001111:	sigmoid = 21'b000000000000000001011;
		14'b10011111010000:	sigmoid = 21'b000000000000000001011;
		14'b10011111010001:	sigmoid = 21'b000000000000000001011;
		14'b10011111010010:	sigmoid = 21'b000000000000000001011;
		14'b10011111010011:	sigmoid = 21'b000000000000000001011;
		14'b10011111010100:	sigmoid = 21'b000000000000000001011;
		14'b10011111010101:	sigmoid = 21'b000000000000000001011;
		14'b10011111010110:	sigmoid = 21'b000000000000000001011;
		14'b10011111010111:	sigmoid = 21'b000000000000000001011;
		14'b10011111011000:	sigmoid = 21'b000000000000000001011;
		14'b10011111011001:	sigmoid = 21'b000000000000000001011;
		14'b10011111011010:	sigmoid = 21'b000000000000000001011;
		14'b10011111011011:	sigmoid = 21'b000000000000000001011;
		14'b10011111011100:	sigmoid = 21'b000000000000000001100;
		14'b10011111011101:	sigmoid = 21'b000000000000000001100;
		14'b10011111011110:	sigmoid = 21'b000000000000000001100;
		14'b10011111011111:	sigmoid = 21'b000000000000000001100;
		14'b10011111100000:	sigmoid = 21'b000000000000000001100;
		14'b10011111100001:	sigmoid = 21'b000000000000000001100;
		14'b10011111100010:	sigmoid = 21'b000000000000000001100;
		14'b10011111100011:	sigmoid = 21'b000000000000000001100;
		14'b10011111100100:	sigmoid = 21'b000000000000000001100;
		14'b10011111100101:	sigmoid = 21'b000000000000000001100;
		14'b10011111100110:	sigmoid = 21'b000000000000000001100;
		14'b10011111100111:	sigmoid = 21'b000000000000000001100;
		14'b10011111101000:	sigmoid = 21'b000000000000000001100;
		14'b10011111101001:	sigmoid = 21'b000000000000000001100;
		14'b10011111101010:	sigmoid = 21'b000000000000000001100;
		14'b10011111101011:	sigmoid = 21'b000000000000000001100;
		14'b10011111101100:	sigmoid = 21'b000000000000000001100;
		14'b10011111101101:	sigmoid = 21'b000000000000000001100;
		14'b10011111101110:	sigmoid = 21'b000000000000000001100;
		14'b10011111101111:	sigmoid = 21'b000000000000000001100;
		14'b10011111110000:	sigmoid = 21'b000000000000000001100;
		14'b10011111110001:	sigmoid = 21'b000000000000000001100;
		14'b10011111110010:	sigmoid = 21'b000000000000000001100;
		14'b10011111110011:	sigmoid = 21'b000000000000000001100;
		14'b10011111110100:	sigmoid = 21'b000000000000000001100;
		14'b10011111110101:	sigmoid = 21'b000000000000000001100;
		14'b10011111110110:	sigmoid = 21'b000000000000000001100;
		14'b10011111110111:	sigmoid = 21'b000000000000000001100;
		14'b10011111111000:	sigmoid = 21'b000000000000000001100;
		14'b10011111111001:	sigmoid = 21'b000000000000000001100;
		14'b10011111111010:	sigmoid = 21'b000000000000000001100;
		14'b10011111111011:	sigmoid = 21'b000000000000000001100;
		14'b10011111111100:	sigmoid = 21'b000000000000000001100;
		14'b10011111111101:	sigmoid = 21'b000000000000000001100;
		14'b10011111111110:	sigmoid = 21'b000000000000000001100;
		14'b10011111111111:	sigmoid = 21'b000000000000000001100;
		14'b10100000000000:	sigmoid = 21'b000000000000000001100;
		14'b10100000000001:	sigmoid = 21'b000000000000000001100;
		14'b10100000000010:	sigmoid = 21'b000000000000000001100;
		14'b10100000000011:	sigmoid = 21'b000000000000000001100;
		14'b10100000000100:	sigmoid = 21'b000000000000000001100;
		14'b10100000000101:	sigmoid = 21'b000000000000000001101;
		14'b10100000000110:	sigmoid = 21'b000000000000000001101;
		14'b10100000000111:	sigmoid = 21'b000000000000000001101;
		14'b10100000001000:	sigmoid = 21'b000000000000000001101;
		14'b10100000001001:	sigmoid = 21'b000000000000000001101;
		14'b10100000001010:	sigmoid = 21'b000000000000000001101;
		14'b10100000001011:	sigmoid = 21'b000000000000000001101;
		14'b10100000001100:	sigmoid = 21'b000000000000000001101;
		14'b10100000001101:	sigmoid = 21'b000000000000000001101;
		14'b10100000001110:	sigmoid = 21'b000000000000000001101;
		14'b10100000001111:	sigmoid = 21'b000000000000000001101;
		14'b10100000010000:	sigmoid = 21'b000000000000000001101;
		14'b10100000010001:	sigmoid = 21'b000000000000000001101;
		14'b10100000010010:	sigmoid = 21'b000000000000000001101;
		14'b10100000010011:	sigmoid = 21'b000000000000000001101;
		14'b10100000010100:	sigmoid = 21'b000000000000000001101;
		14'b10100000010101:	sigmoid = 21'b000000000000000001101;
		14'b10100000010110:	sigmoid = 21'b000000000000000001101;
		14'b10100000010111:	sigmoid = 21'b000000000000000001101;
		14'b10100000011000:	sigmoid = 21'b000000000000000001101;
		14'b10100000011001:	sigmoid = 21'b000000000000000001101;
		14'b10100000011010:	sigmoid = 21'b000000000000000001101;
		14'b10100000011011:	sigmoid = 21'b000000000000000001101;
		14'b10100000011100:	sigmoid = 21'b000000000000000001101;
		14'b10100000011101:	sigmoid = 21'b000000000000000001101;
		14'b10100000011110:	sigmoid = 21'b000000000000000001101;
		14'b10100000011111:	sigmoid = 21'b000000000000000001101;
		14'b10100000100000:	sigmoid = 21'b000000000000000001101;
		14'b10100000100001:	sigmoid = 21'b000000000000000001101;
		14'b10100000100010:	sigmoid = 21'b000000000000000001101;
		14'b10100000100011:	sigmoid = 21'b000000000000000001101;
		14'b10100000100100:	sigmoid = 21'b000000000000000001101;
		14'b10100000100101:	sigmoid = 21'b000000000000000001101;
		14'b10100000100110:	sigmoid = 21'b000000000000000001101;
		14'b10100000100111:	sigmoid = 21'b000000000000000001101;
		14'b10100000101000:	sigmoid = 21'b000000000000000001101;
		14'b10100000101001:	sigmoid = 21'b000000000000000001101;
		14'b10100000101010:	sigmoid = 21'b000000000000000001101;
		14'b10100000101011:	sigmoid = 21'b000000000000000001110;
		14'b10100000101100:	sigmoid = 21'b000000000000000001110;
		14'b10100000101101:	sigmoid = 21'b000000000000000001110;
		14'b10100000101110:	sigmoid = 21'b000000000000000001110;
		14'b10100000101111:	sigmoid = 21'b000000000000000001110;
		14'b10100000110000:	sigmoid = 21'b000000000000000001110;
		14'b10100000110001:	sigmoid = 21'b000000000000000001110;
		14'b10100000110010:	sigmoid = 21'b000000000000000001110;
		14'b10100000110011:	sigmoid = 21'b000000000000000001110;
		14'b10100000110100:	sigmoid = 21'b000000000000000001110;
		14'b10100000110101:	sigmoid = 21'b000000000000000001110;
		14'b10100000110110:	sigmoid = 21'b000000000000000001110;
		14'b10100000110111:	sigmoid = 21'b000000000000000001110;
		14'b10100000111000:	sigmoid = 21'b000000000000000001110;
		14'b10100000111001:	sigmoid = 21'b000000000000000001110;
		14'b10100000111010:	sigmoid = 21'b000000000000000001110;
		14'b10100000111011:	sigmoid = 21'b000000000000000001110;
		14'b10100000111100:	sigmoid = 21'b000000000000000001110;
		14'b10100000111101:	sigmoid = 21'b000000000000000001110;
		14'b10100000111110:	sigmoid = 21'b000000000000000001110;
		14'b10100000111111:	sigmoid = 21'b000000000000000001110;
		14'b10100001000000:	sigmoid = 21'b000000000000000001110;
		14'b10100001000001:	sigmoid = 21'b000000000000000001110;
		14'b10100001000010:	sigmoid = 21'b000000000000000001110;
		14'b10100001000011:	sigmoid = 21'b000000000000000001110;
		14'b10100001000100:	sigmoid = 21'b000000000000000001110;
		14'b10100001000101:	sigmoid = 21'b000000000000000001110;
		14'b10100001000110:	sigmoid = 21'b000000000000000001110;
		14'b10100001000111:	sigmoid = 21'b000000000000000001110;
		14'b10100001001000:	sigmoid = 21'b000000000000000001110;
		14'b10100001001001:	sigmoid = 21'b000000000000000001110;
		14'b10100001001010:	sigmoid = 21'b000000000000000001110;
		14'b10100001001011:	sigmoid = 21'b000000000000000001110;
		14'b10100001001100:	sigmoid = 21'b000000000000000001110;
		14'b10100001001101:	sigmoid = 21'b000000000000000001110;
		14'b10100001001110:	sigmoid = 21'b000000000000000001111;
		14'b10100001001111:	sigmoid = 21'b000000000000000001111;
		14'b10100001010000:	sigmoid = 21'b000000000000000001111;
		14'b10100001010001:	sigmoid = 21'b000000000000000001111;
		14'b10100001010010:	sigmoid = 21'b000000000000000001111;
		14'b10100001010011:	sigmoid = 21'b000000000000000001111;
		14'b10100001010100:	sigmoid = 21'b000000000000000001111;
		14'b10100001010101:	sigmoid = 21'b000000000000000001111;
		14'b10100001010110:	sigmoid = 21'b000000000000000001111;
		14'b10100001010111:	sigmoid = 21'b000000000000000001111;
		14'b10100001011000:	sigmoid = 21'b000000000000000001111;
		14'b10100001011001:	sigmoid = 21'b000000000000000001111;
		14'b10100001011010:	sigmoid = 21'b000000000000000001111;
		14'b10100001011011:	sigmoid = 21'b000000000000000001111;
		14'b10100001011100:	sigmoid = 21'b000000000000000001111;
		14'b10100001011101:	sigmoid = 21'b000000000000000001111;
		14'b10100001011110:	sigmoid = 21'b000000000000000001111;
		14'b10100001011111:	sigmoid = 21'b000000000000000001111;
		14'b10100001100000:	sigmoid = 21'b000000000000000001111;
		14'b10100001100001:	sigmoid = 21'b000000000000000001111;
		14'b10100001100010:	sigmoid = 21'b000000000000000001111;
		14'b10100001100011:	sigmoid = 21'b000000000000000001111;
		14'b10100001100100:	sigmoid = 21'b000000000000000001111;
		14'b10100001100101:	sigmoid = 21'b000000000000000001111;
		14'b10100001100110:	sigmoid = 21'b000000000000000001111;
		14'b10100001100111:	sigmoid = 21'b000000000000000001111;
		14'b10100001101000:	sigmoid = 21'b000000000000000001111;
		14'b10100001101001:	sigmoid = 21'b000000000000000001111;
		14'b10100001101010:	sigmoid = 21'b000000000000000001111;
		14'b10100001101011:	sigmoid = 21'b000000000000000001111;
		14'b10100001101100:	sigmoid = 21'b000000000000000001111;
		14'b10100001101101:	sigmoid = 21'b000000000000000001111;
		14'b10100001101110:	sigmoid = 21'b000000000000000001111;
		14'b10100001101111:	sigmoid = 21'b000000000000000010000;
		14'b10100001110000:	sigmoid = 21'b000000000000000010000;
		14'b10100001110001:	sigmoid = 21'b000000000000000010000;
		14'b10100001110010:	sigmoid = 21'b000000000000000010000;
		14'b10100001110011:	sigmoid = 21'b000000000000000010000;
		14'b10100001110100:	sigmoid = 21'b000000000000000010000;
		14'b10100001110101:	sigmoid = 21'b000000000000000010000;
		14'b10100001110110:	sigmoid = 21'b000000000000000010000;
		14'b10100001110111:	sigmoid = 21'b000000000000000010000;
		14'b10100001111000:	sigmoid = 21'b000000000000000010000;
		14'b10100001111001:	sigmoid = 21'b000000000000000010000;
		14'b10100001111010:	sigmoid = 21'b000000000000000010000;
		14'b10100001111011:	sigmoid = 21'b000000000000000010000;
		14'b10100001111100:	sigmoid = 21'b000000000000000010000;
		14'b10100001111101:	sigmoid = 21'b000000000000000010000;
		14'b10100001111110:	sigmoid = 21'b000000000000000010000;
		14'b10100001111111:	sigmoid = 21'b000000000000000010000;
		14'b10100010000000:	sigmoid = 21'b000000000000000010000;
		14'b10100010000001:	sigmoid = 21'b000000000000000010000;
		14'b10100010000010:	sigmoid = 21'b000000000000000010000;
		14'b10100010000011:	sigmoid = 21'b000000000000000010000;
		14'b10100010000100:	sigmoid = 21'b000000000000000010000;
		14'b10100010000101:	sigmoid = 21'b000000000000000010000;
		14'b10100010000110:	sigmoid = 21'b000000000000000010000;
		14'b10100010000111:	sigmoid = 21'b000000000000000010000;
		14'b10100010001000:	sigmoid = 21'b000000000000000010000;
		14'b10100010001001:	sigmoid = 21'b000000000000000010000;
		14'b10100010001010:	sigmoid = 21'b000000000000000010000;
		14'b10100010001011:	sigmoid = 21'b000000000000000010000;
		14'b10100010001100:	sigmoid = 21'b000000000000000010000;
		14'b10100010001101:	sigmoid = 21'b000000000000000010000;
		14'b10100010001110:	sigmoid = 21'b000000000000000010001;
		14'b10100010001111:	sigmoid = 21'b000000000000000010001;
		14'b10100010010000:	sigmoid = 21'b000000000000000010001;
		14'b10100010010001:	sigmoid = 21'b000000000000000010001;
		14'b10100010010010:	sigmoid = 21'b000000000000000010001;
		14'b10100010010011:	sigmoid = 21'b000000000000000010001;
		14'b10100010010100:	sigmoid = 21'b000000000000000010001;
		14'b10100010010101:	sigmoid = 21'b000000000000000010001;
		14'b10100010010110:	sigmoid = 21'b000000000000000010001;
		14'b10100010010111:	sigmoid = 21'b000000000000000010001;
		14'b10100010011000:	sigmoid = 21'b000000000000000010001;
		14'b10100010011001:	sigmoid = 21'b000000000000000010001;
		14'b10100010011010:	sigmoid = 21'b000000000000000010001;
		14'b10100010011011:	sigmoid = 21'b000000000000000010001;
		14'b10100010011100:	sigmoid = 21'b000000000000000010001;
		14'b10100010011101:	sigmoid = 21'b000000000000000010001;
		14'b10100010011110:	sigmoid = 21'b000000000000000010001;
		14'b10100010011111:	sigmoid = 21'b000000000000000010001;
		14'b10100010100000:	sigmoid = 21'b000000000000000010001;
		14'b10100010100001:	sigmoid = 21'b000000000000000010001;
		14'b10100010100010:	sigmoid = 21'b000000000000000010001;
		14'b10100010100011:	sigmoid = 21'b000000000000000010001;
		14'b10100010100100:	sigmoid = 21'b000000000000000010001;
		14'b10100010100101:	sigmoid = 21'b000000000000000010001;
		14'b10100010100110:	sigmoid = 21'b000000000000000010001;
		14'b10100010100111:	sigmoid = 21'b000000000000000010001;
		14'b10100010101000:	sigmoid = 21'b000000000000000010001;
		14'b10100010101001:	sigmoid = 21'b000000000000000010001;
		14'b10100010101010:	sigmoid = 21'b000000000000000010001;
		14'b10100010101011:	sigmoid = 21'b000000000000000010001;
		14'b10100010101100:	sigmoid = 21'b000000000000000010010;
		14'b10100010101101:	sigmoid = 21'b000000000000000010010;
		14'b10100010101110:	sigmoid = 21'b000000000000000010010;
		14'b10100010101111:	sigmoid = 21'b000000000000000010010;
		14'b10100010110000:	sigmoid = 21'b000000000000000010010;
		14'b10100010110001:	sigmoid = 21'b000000000000000010010;
		14'b10100010110010:	sigmoid = 21'b000000000000000010010;
		14'b10100010110011:	sigmoid = 21'b000000000000000010010;
		14'b10100010110100:	sigmoid = 21'b000000000000000010010;
		14'b10100010110101:	sigmoid = 21'b000000000000000010010;
		14'b10100010110110:	sigmoid = 21'b000000000000000010010;
		14'b10100010110111:	sigmoid = 21'b000000000000000010010;
		14'b10100010111000:	sigmoid = 21'b000000000000000010010;
		14'b10100010111001:	sigmoid = 21'b000000000000000010010;
		14'b10100010111010:	sigmoid = 21'b000000000000000010010;
		14'b10100010111011:	sigmoid = 21'b000000000000000010010;
		14'b10100010111100:	sigmoid = 21'b000000000000000010010;
		14'b10100010111101:	sigmoid = 21'b000000000000000010010;
		14'b10100010111110:	sigmoid = 21'b000000000000000010010;
		14'b10100010111111:	sigmoid = 21'b000000000000000010010;
		14'b10100011000000:	sigmoid = 21'b000000000000000010010;
		14'b10100011000001:	sigmoid = 21'b000000000000000010010;
		14'b10100011000010:	sigmoid = 21'b000000000000000010010;
		14'b10100011000011:	sigmoid = 21'b000000000000000010010;
		14'b10100011000100:	sigmoid = 21'b000000000000000010010;
		14'b10100011000101:	sigmoid = 21'b000000000000000010010;
		14'b10100011000110:	sigmoid = 21'b000000000000000010010;
		14'b10100011000111:	sigmoid = 21'b000000000000000010011;
		14'b10100011001000:	sigmoid = 21'b000000000000000010011;
		14'b10100011001001:	sigmoid = 21'b000000000000000010011;
		14'b10100011001010:	sigmoid = 21'b000000000000000010011;
		14'b10100011001011:	sigmoid = 21'b000000000000000010011;
		14'b10100011001100:	sigmoid = 21'b000000000000000010011;
		14'b10100011001101:	sigmoid = 21'b000000000000000010011;
		14'b10100011001110:	sigmoid = 21'b000000000000000010011;
		14'b10100011001111:	sigmoid = 21'b000000000000000010011;
		14'b10100011010000:	sigmoid = 21'b000000000000000010011;
		14'b10100011010001:	sigmoid = 21'b000000000000000010011;
		14'b10100011010010:	sigmoid = 21'b000000000000000010011;
		14'b10100011010011:	sigmoid = 21'b000000000000000010011;
		14'b10100011010100:	sigmoid = 21'b000000000000000010011;
		14'b10100011010101:	sigmoid = 21'b000000000000000010011;
		14'b10100011010110:	sigmoid = 21'b000000000000000010011;
		14'b10100011010111:	sigmoid = 21'b000000000000000010011;
		14'b10100011011000:	sigmoid = 21'b000000000000000010011;
		14'b10100011011001:	sigmoid = 21'b000000000000000010011;
		14'b10100011011010:	sigmoid = 21'b000000000000000010011;
		14'b10100011011011:	sigmoid = 21'b000000000000000010011;
		14'b10100011011100:	sigmoid = 21'b000000000000000010011;
		14'b10100011011101:	sigmoid = 21'b000000000000000010011;
		14'b10100011011110:	sigmoid = 21'b000000000000000010011;
		14'b10100011011111:	sigmoid = 21'b000000000000000010011;
		14'b10100011100000:	sigmoid = 21'b000000000000000010011;
		14'b10100011100001:	sigmoid = 21'b000000000000000010011;
		14'b10100011100010:	sigmoid = 21'b000000000000000010100;
		14'b10100011100011:	sigmoid = 21'b000000000000000010100;
		14'b10100011100100:	sigmoid = 21'b000000000000000010100;
		14'b10100011100101:	sigmoid = 21'b000000000000000010100;
		14'b10100011100110:	sigmoid = 21'b000000000000000010100;
		14'b10100011100111:	sigmoid = 21'b000000000000000010100;
		14'b10100011101000:	sigmoid = 21'b000000000000000010100;
		14'b10100011101001:	sigmoid = 21'b000000000000000010100;
		14'b10100011101010:	sigmoid = 21'b000000000000000010100;
		14'b10100011101011:	sigmoid = 21'b000000000000000010100;
		14'b10100011101100:	sigmoid = 21'b000000000000000010100;
		14'b10100011101101:	sigmoid = 21'b000000000000000010100;
		14'b10100011101110:	sigmoid = 21'b000000000000000010100;
		14'b10100011101111:	sigmoid = 21'b000000000000000010100;
		14'b10100011110000:	sigmoid = 21'b000000000000000010100;
		14'b10100011110001:	sigmoid = 21'b000000000000000010100;
		14'b10100011110010:	sigmoid = 21'b000000000000000010100;
		14'b10100011110011:	sigmoid = 21'b000000000000000010100;
		14'b10100011110100:	sigmoid = 21'b000000000000000010100;
		14'b10100011110101:	sigmoid = 21'b000000000000000010100;
		14'b10100011110110:	sigmoid = 21'b000000000000000010100;
		14'b10100011110111:	sigmoid = 21'b000000000000000010100;
		14'b10100011111000:	sigmoid = 21'b000000000000000010100;
		14'b10100011111001:	sigmoid = 21'b000000000000000010100;
		14'b10100011111010:	sigmoid = 21'b000000000000000010100;
		14'b10100011111011:	sigmoid = 21'b000000000000000010101;
		14'b10100011111100:	sigmoid = 21'b000000000000000010101;
		14'b10100011111101:	sigmoid = 21'b000000000000000010101;
		14'b10100011111110:	sigmoid = 21'b000000000000000010101;
		14'b10100011111111:	sigmoid = 21'b000000000000000010101;
		14'b10100100000000:	sigmoid = 21'b000000000000000010101;
		14'b10100100000001:	sigmoid = 21'b000000000000000010101;
		14'b10100100000010:	sigmoid = 21'b000000000000000010101;
		14'b10100100000011:	sigmoid = 21'b000000000000000010101;
		14'b10100100000100:	sigmoid = 21'b000000000000000010101;
		14'b10100100000101:	sigmoid = 21'b000000000000000010101;
		14'b10100100000110:	sigmoid = 21'b000000000000000010101;
		14'b10100100000111:	sigmoid = 21'b000000000000000010101;
		14'b10100100001000:	sigmoid = 21'b000000000000000010101;
		14'b10100100001001:	sigmoid = 21'b000000000000000010101;
		14'b10100100001010:	sigmoid = 21'b000000000000000010101;
		14'b10100100001011:	sigmoid = 21'b000000000000000010101;
		14'b10100100001100:	sigmoid = 21'b000000000000000010101;
		14'b10100100001101:	sigmoid = 21'b000000000000000010101;
		14'b10100100001110:	sigmoid = 21'b000000000000000010101;
		14'b10100100001111:	sigmoid = 21'b000000000000000010101;
		14'b10100100010000:	sigmoid = 21'b000000000000000010101;
		14'b10100100010001:	sigmoid = 21'b000000000000000010101;
		14'b10100100010010:	sigmoid = 21'b000000000000000010110;
		14'b10100100010011:	sigmoid = 21'b000000000000000010110;
		14'b10100100010100:	sigmoid = 21'b000000000000000010110;
		14'b10100100010101:	sigmoid = 21'b000000000000000010110;
		14'b10100100010110:	sigmoid = 21'b000000000000000010110;
		14'b10100100010111:	sigmoid = 21'b000000000000000010110;
		14'b10100100011000:	sigmoid = 21'b000000000000000010110;
		14'b10100100011001:	sigmoid = 21'b000000000000000010110;
		14'b10100100011010:	sigmoid = 21'b000000000000000010110;
		14'b10100100011011:	sigmoid = 21'b000000000000000010110;
		14'b10100100011100:	sigmoid = 21'b000000000000000010110;
		14'b10100100011101:	sigmoid = 21'b000000000000000010110;
		14'b10100100011110:	sigmoid = 21'b000000000000000010110;
		14'b10100100011111:	sigmoid = 21'b000000000000000010110;
		14'b10100100100000:	sigmoid = 21'b000000000000000010110;
		14'b10100100100001:	sigmoid = 21'b000000000000000010110;
		14'b10100100100010:	sigmoid = 21'b000000000000000010110;
		14'b10100100100011:	sigmoid = 21'b000000000000000010110;
		14'b10100100100100:	sigmoid = 21'b000000000000000010110;
		14'b10100100100101:	sigmoid = 21'b000000000000000010110;
		14'b10100100100110:	sigmoid = 21'b000000000000000010110;
		14'b10100100100111:	sigmoid = 21'b000000000000000010110;
		14'b10100100101000:	sigmoid = 21'b000000000000000010110;
		14'b10100100101001:	sigmoid = 21'b000000000000000010111;
		14'b10100100101010:	sigmoid = 21'b000000000000000010111;
		14'b10100100101011:	sigmoid = 21'b000000000000000010111;
		14'b10100100101100:	sigmoid = 21'b000000000000000010111;
		14'b10100100101101:	sigmoid = 21'b000000000000000010111;
		14'b10100100101110:	sigmoid = 21'b000000000000000010111;
		14'b10100100101111:	sigmoid = 21'b000000000000000010111;
		14'b10100100110000:	sigmoid = 21'b000000000000000010111;
		14'b10100100110001:	sigmoid = 21'b000000000000000010111;
		14'b10100100110010:	sigmoid = 21'b000000000000000010111;
		14'b10100100110011:	sigmoid = 21'b000000000000000010111;
		14'b10100100110100:	sigmoid = 21'b000000000000000010111;
		14'b10100100110101:	sigmoid = 21'b000000000000000010111;
		14'b10100100110110:	sigmoid = 21'b000000000000000010111;
		14'b10100100110111:	sigmoid = 21'b000000000000000010111;
		14'b10100100111000:	sigmoid = 21'b000000000000000010111;
		14'b10100100111001:	sigmoid = 21'b000000000000000010111;
		14'b10100100111010:	sigmoid = 21'b000000000000000010111;
		14'b10100100111011:	sigmoid = 21'b000000000000000010111;
		14'b10100100111100:	sigmoid = 21'b000000000000000010111;
		14'b10100100111101:	sigmoid = 21'b000000000000000010111;
		14'b10100100111110:	sigmoid = 21'b000000000000000010111;
		14'b10100100111111:	sigmoid = 21'b000000000000000011000;
		14'b10100101000000:	sigmoid = 21'b000000000000000011000;
		14'b10100101000001:	sigmoid = 21'b000000000000000011000;
		14'b10100101000010:	sigmoid = 21'b000000000000000011000;
		14'b10100101000011:	sigmoid = 21'b000000000000000011000;
		14'b10100101000100:	sigmoid = 21'b000000000000000011000;
		14'b10100101000101:	sigmoid = 21'b000000000000000011000;
		14'b10100101000110:	sigmoid = 21'b000000000000000011000;
		14'b10100101000111:	sigmoid = 21'b000000000000000011000;
		14'b10100101001000:	sigmoid = 21'b000000000000000011000;
		14'b10100101001001:	sigmoid = 21'b000000000000000011000;
		14'b10100101001010:	sigmoid = 21'b000000000000000011000;
		14'b10100101001011:	sigmoid = 21'b000000000000000011000;
		14'b10100101001100:	sigmoid = 21'b000000000000000011000;
		14'b10100101001101:	sigmoid = 21'b000000000000000011000;
		14'b10100101001110:	sigmoid = 21'b000000000000000011000;
		14'b10100101001111:	sigmoid = 21'b000000000000000011000;
		14'b10100101010000:	sigmoid = 21'b000000000000000011000;
		14'b10100101010001:	sigmoid = 21'b000000000000000011000;
		14'b10100101010010:	sigmoid = 21'b000000000000000011000;
		14'b10100101010011:	sigmoid = 21'b000000000000000011000;
		14'b10100101010100:	sigmoid = 21'b000000000000000011001;
		14'b10100101010101:	sigmoid = 21'b000000000000000011001;
		14'b10100101010110:	sigmoid = 21'b000000000000000011001;
		14'b10100101010111:	sigmoid = 21'b000000000000000011001;
		14'b10100101011000:	sigmoid = 21'b000000000000000011001;
		14'b10100101011001:	sigmoid = 21'b000000000000000011001;
		14'b10100101011010:	sigmoid = 21'b000000000000000011001;
		14'b10100101011011:	sigmoid = 21'b000000000000000011001;
		14'b10100101011100:	sigmoid = 21'b000000000000000011001;
		14'b10100101011101:	sigmoid = 21'b000000000000000011001;
		14'b10100101011110:	sigmoid = 21'b000000000000000011001;
		14'b10100101011111:	sigmoid = 21'b000000000000000011001;
		14'b10100101100000:	sigmoid = 21'b000000000000000011001;
		14'b10100101100001:	sigmoid = 21'b000000000000000011001;
		14'b10100101100010:	sigmoid = 21'b000000000000000011001;
		14'b10100101100011:	sigmoid = 21'b000000000000000011001;
		14'b10100101100100:	sigmoid = 21'b000000000000000011001;
		14'b10100101100101:	sigmoid = 21'b000000000000000011001;
		14'b10100101100110:	sigmoid = 21'b000000000000000011001;
		14'b10100101100111:	sigmoid = 21'b000000000000000011001;
		14'b10100101101000:	sigmoid = 21'b000000000000000011010;
		14'b10100101101001:	sigmoid = 21'b000000000000000011010;
		14'b10100101101010:	sigmoid = 21'b000000000000000011010;
		14'b10100101101011:	sigmoid = 21'b000000000000000011010;
		14'b10100101101100:	sigmoid = 21'b000000000000000011010;
		14'b10100101101101:	sigmoid = 21'b000000000000000011010;
		14'b10100101101110:	sigmoid = 21'b000000000000000011010;
		14'b10100101101111:	sigmoid = 21'b000000000000000011010;
		14'b10100101110000:	sigmoid = 21'b000000000000000011010;
		14'b10100101110001:	sigmoid = 21'b000000000000000011010;
		14'b10100101110010:	sigmoid = 21'b000000000000000011010;
		14'b10100101110011:	sigmoid = 21'b000000000000000011010;
		14'b10100101110100:	sigmoid = 21'b000000000000000011010;
		14'b10100101110101:	sigmoid = 21'b000000000000000011010;
		14'b10100101110110:	sigmoid = 21'b000000000000000011010;
		14'b10100101110111:	sigmoid = 21'b000000000000000011010;
		14'b10100101111000:	sigmoid = 21'b000000000000000011010;
		14'b10100101111001:	sigmoid = 21'b000000000000000011010;
		14'b10100101111010:	sigmoid = 21'b000000000000000011010;
		14'b10100101111011:	sigmoid = 21'b000000000000000011011;
		14'b10100101111100:	sigmoid = 21'b000000000000000011011;
		14'b10100101111101:	sigmoid = 21'b000000000000000011011;
		14'b10100101111110:	sigmoid = 21'b000000000000000011011;
		14'b10100101111111:	sigmoid = 21'b000000000000000011011;
		14'b10100110000000:	sigmoid = 21'b000000000000000011011;
		14'b10100110000001:	sigmoid = 21'b000000000000000011011;
		14'b10100110000010:	sigmoid = 21'b000000000000000011011;
		14'b10100110000011:	sigmoid = 21'b000000000000000011011;
		14'b10100110000100:	sigmoid = 21'b000000000000000011011;
		14'b10100110000101:	sigmoid = 21'b000000000000000011011;
		14'b10100110000110:	sigmoid = 21'b000000000000000011011;
		14'b10100110000111:	sigmoid = 21'b000000000000000011011;
		14'b10100110001000:	sigmoid = 21'b000000000000000011011;
		14'b10100110001001:	sigmoid = 21'b000000000000000011011;
		14'b10100110001010:	sigmoid = 21'b000000000000000011011;
		14'b10100110001011:	sigmoid = 21'b000000000000000011011;
		14'b10100110001100:	sigmoid = 21'b000000000000000011011;
		14'b10100110001101:	sigmoid = 21'b000000000000000011011;
		14'b10100110001110:	sigmoid = 21'b000000000000000011100;
		14'b10100110001111:	sigmoid = 21'b000000000000000011100;
		14'b10100110010000:	sigmoid = 21'b000000000000000011100;
		14'b10100110010001:	sigmoid = 21'b000000000000000011100;
		14'b10100110010010:	sigmoid = 21'b000000000000000011100;
		14'b10100110010011:	sigmoid = 21'b000000000000000011100;
		14'b10100110010100:	sigmoid = 21'b000000000000000011100;
		14'b10100110010101:	sigmoid = 21'b000000000000000011100;
		14'b10100110010110:	sigmoid = 21'b000000000000000011100;
		14'b10100110010111:	sigmoid = 21'b000000000000000011100;
		14'b10100110011000:	sigmoid = 21'b000000000000000011100;
		14'b10100110011001:	sigmoid = 21'b000000000000000011100;
		14'b10100110011010:	sigmoid = 21'b000000000000000011100;
		14'b10100110011011:	sigmoid = 21'b000000000000000011100;
		14'b10100110011100:	sigmoid = 21'b000000000000000011100;
		14'b10100110011101:	sigmoid = 21'b000000000000000011100;
		14'b10100110011110:	sigmoid = 21'b000000000000000011100;
		14'b10100110011111:	sigmoid = 21'b000000000000000011100;
		14'b10100110100000:	sigmoid = 21'b000000000000000011101;
		14'b10100110100001:	sigmoid = 21'b000000000000000011101;
		14'b10100110100010:	sigmoid = 21'b000000000000000011101;
		14'b10100110100011:	sigmoid = 21'b000000000000000011101;
		14'b10100110100100:	sigmoid = 21'b000000000000000011101;
		14'b10100110100101:	sigmoid = 21'b000000000000000011101;
		14'b10100110100110:	sigmoid = 21'b000000000000000011101;
		14'b10100110100111:	sigmoid = 21'b000000000000000011101;
		14'b10100110101000:	sigmoid = 21'b000000000000000011101;
		14'b10100110101001:	sigmoid = 21'b000000000000000011101;
		14'b10100110101010:	sigmoid = 21'b000000000000000011101;
		14'b10100110101011:	sigmoid = 21'b000000000000000011101;
		14'b10100110101100:	sigmoid = 21'b000000000000000011101;
		14'b10100110101101:	sigmoid = 21'b000000000000000011101;
		14'b10100110101110:	sigmoid = 21'b000000000000000011101;
		14'b10100110101111:	sigmoid = 21'b000000000000000011101;
		14'b10100110110000:	sigmoid = 21'b000000000000000011101;
		14'b10100110110001:	sigmoid = 21'b000000000000000011110;
		14'b10100110110010:	sigmoid = 21'b000000000000000011110;
		14'b10100110110011:	sigmoid = 21'b000000000000000011110;
		14'b10100110110100:	sigmoid = 21'b000000000000000011110;
		14'b10100110110101:	sigmoid = 21'b000000000000000011110;
		14'b10100110110110:	sigmoid = 21'b000000000000000011110;
		14'b10100110110111:	sigmoid = 21'b000000000000000011110;
		14'b10100110111000:	sigmoid = 21'b000000000000000011110;
		14'b10100110111001:	sigmoid = 21'b000000000000000011110;
		14'b10100110111010:	sigmoid = 21'b000000000000000011110;
		14'b10100110111011:	sigmoid = 21'b000000000000000011110;
		14'b10100110111100:	sigmoid = 21'b000000000000000011110;
		14'b10100110111101:	sigmoid = 21'b000000000000000011110;
		14'b10100110111110:	sigmoid = 21'b000000000000000011110;
		14'b10100110111111:	sigmoid = 21'b000000000000000011110;
		14'b10100111000000:	sigmoid = 21'b000000000000000011110;
		14'b10100111000001:	sigmoid = 21'b000000000000000011110;
		14'b10100111000010:	sigmoid = 21'b000000000000000011111;
		14'b10100111000011:	sigmoid = 21'b000000000000000011111;
		14'b10100111000100:	sigmoid = 21'b000000000000000011111;
		14'b10100111000101:	sigmoid = 21'b000000000000000011111;
		14'b10100111000110:	sigmoid = 21'b000000000000000011111;
		14'b10100111000111:	sigmoid = 21'b000000000000000011111;
		14'b10100111001000:	sigmoid = 21'b000000000000000011111;
		14'b10100111001001:	sigmoid = 21'b000000000000000011111;
		14'b10100111001010:	sigmoid = 21'b000000000000000011111;
		14'b10100111001011:	sigmoid = 21'b000000000000000011111;
		14'b10100111001100:	sigmoid = 21'b000000000000000011111;
		14'b10100111001101:	sigmoid = 21'b000000000000000011111;
		14'b10100111001110:	sigmoid = 21'b000000000000000011111;
		14'b10100111001111:	sigmoid = 21'b000000000000000011111;
		14'b10100111010000:	sigmoid = 21'b000000000000000011111;
		14'b10100111010001:	sigmoid = 21'b000000000000000011111;
		14'b10100111010010:	sigmoid = 21'b000000000000000100000;
		14'b10100111010011:	sigmoid = 21'b000000000000000100000;
		14'b10100111010100:	sigmoid = 21'b000000000000000100000;
		14'b10100111010101:	sigmoid = 21'b000000000000000100000;
		14'b10100111010110:	sigmoid = 21'b000000000000000100000;
		14'b10100111010111:	sigmoid = 21'b000000000000000100000;
		14'b10100111011000:	sigmoid = 21'b000000000000000100000;
		14'b10100111011001:	sigmoid = 21'b000000000000000100000;
		14'b10100111011010:	sigmoid = 21'b000000000000000100000;
		14'b10100111011011:	sigmoid = 21'b000000000000000100000;
		14'b10100111011100:	sigmoid = 21'b000000000000000100000;
		14'b10100111011101:	sigmoid = 21'b000000000000000100000;
		14'b10100111011110:	sigmoid = 21'b000000000000000100000;
		14'b10100111011111:	sigmoid = 21'b000000000000000100000;
		14'b10100111100000:	sigmoid = 21'b000000000000000100000;
		14'b10100111100001:	sigmoid = 21'b000000000000000100000;
		14'b10100111100010:	sigmoid = 21'b000000000000000100001;
		14'b10100111100011:	sigmoid = 21'b000000000000000100001;
		14'b10100111100100:	sigmoid = 21'b000000000000000100001;
		14'b10100111100101:	sigmoid = 21'b000000000000000100001;
		14'b10100111100110:	sigmoid = 21'b000000000000000100001;
		14'b10100111100111:	sigmoid = 21'b000000000000000100001;
		14'b10100111101000:	sigmoid = 21'b000000000000000100001;
		14'b10100111101001:	sigmoid = 21'b000000000000000100001;
		14'b10100111101010:	sigmoid = 21'b000000000000000100001;
		14'b10100111101011:	sigmoid = 21'b000000000000000100001;
		14'b10100111101100:	sigmoid = 21'b000000000000000100001;
		14'b10100111101101:	sigmoid = 21'b000000000000000100001;
		14'b10100111101110:	sigmoid = 21'b000000000000000100001;
		14'b10100111101111:	sigmoid = 21'b000000000000000100001;
		14'b10100111110000:	sigmoid = 21'b000000000000000100001;
		14'b10100111110001:	sigmoid = 21'b000000000000000100010;
		14'b10100111110010:	sigmoid = 21'b000000000000000100010;
		14'b10100111110011:	sigmoid = 21'b000000000000000100010;
		14'b10100111110100:	sigmoid = 21'b000000000000000100010;
		14'b10100111110101:	sigmoid = 21'b000000000000000100010;
		14'b10100111110110:	sigmoid = 21'b000000000000000100010;
		14'b10100111110111:	sigmoid = 21'b000000000000000100010;
		14'b10100111111000:	sigmoid = 21'b000000000000000100010;
		14'b10100111111001:	sigmoid = 21'b000000000000000100010;
		14'b10100111111010:	sigmoid = 21'b000000000000000100010;
		14'b10100111111011:	sigmoid = 21'b000000000000000100010;
		14'b10100111111100:	sigmoid = 21'b000000000000000100010;
		14'b10100111111101:	sigmoid = 21'b000000000000000100010;
		14'b10100111111110:	sigmoid = 21'b000000000000000100010;
		14'b10100111111111:	sigmoid = 21'b000000000000000100010;
		14'b10101000000000:	sigmoid = 21'b000000000000000100011;
		14'b10101000000001:	sigmoid = 21'b000000000000000100011;
		14'b10101000000010:	sigmoid = 21'b000000000000000100011;
		14'b10101000000011:	sigmoid = 21'b000000000000000100011;
		14'b10101000000100:	sigmoid = 21'b000000000000000100011;
		14'b10101000000101:	sigmoid = 21'b000000000000000100011;
		14'b10101000000110:	sigmoid = 21'b000000000000000100011;
		14'b10101000000111:	sigmoid = 21'b000000000000000100011;
		14'b10101000001000:	sigmoid = 21'b000000000000000100011;
		14'b10101000001001:	sigmoid = 21'b000000000000000100011;
		14'b10101000001010:	sigmoid = 21'b000000000000000100011;
		14'b10101000001011:	sigmoid = 21'b000000000000000100011;
		14'b10101000001100:	sigmoid = 21'b000000000000000100011;
		14'b10101000001101:	sigmoid = 21'b000000000000000100011;
		14'b10101000001110:	sigmoid = 21'b000000000000000100011;
		14'b10101000001111:	sigmoid = 21'b000000000000000100100;
		14'b10101000010000:	sigmoid = 21'b000000000000000100100;
		14'b10101000010001:	sigmoid = 21'b000000000000000100100;
		14'b10101000010010:	sigmoid = 21'b000000000000000100100;
		14'b10101000010011:	sigmoid = 21'b000000000000000100100;
		14'b10101000010100:	sigmoid = 21'b000000000000000100100;
		14'b10101000010101:	sigmoid = 21'b000000000000000100100;
		14'b10101000010110:	sigmoid = 21'b000000000000000100100;
		14'b10101000010111:	sigmoid = 21'b000000000000000100100;
		14'b10101000011000:	sigmoid = 21'b000000000000000100100;
		14'b10101000011001:	sigmoid = 21'b000000000000000100100;
		14'b10101000011010:	sigmoid = 21'b000000000000000100100;
		14'b10101000011011:	sigmoid = 21'b000000000000000100100;
		14'b10101000011100:	sigmoid = 21'b000000000000000100100;
		14'b10101000011101:	sigmoid = 21'b000000000000000100101;
		14'b10101000011110:	sigmoid = 21'b000000000000000100101;
		14'b10101000011111:	sigmoid = 21'b000000000000000100101;
		14'b10101000100000:	sigmoid = 21'b000000000000000100101;
		14'b10101000100001:	sigmoid = 21'b000000000000000100101;
		14'b10101000100010:	sigmoid = 21'b000000000000000100101;
		14'b10101000100011:	sigmoid = 21'b000000000000000100101;
		14'b10101000100100:	sigmoid = 21'b000000000000000100101;
		14'b10101000100101:	sigmoid = 21'b000000000000000100101;
		14'b10101000100110:	sigmoid = 21'b000000000000000100101;
		14'b10101000100111:	sigmoid = 21'b000000000000000100101;
		14'b10101000101000:	sigmoid = 21'b000000000000000100101;
		14'b10101000101001:	sigmoid = 21'b000000000000000100101;
		14'b10101000101010:	sigmoid = 21'b000000000000000100110;
		14'b10101000101011:	sigmoid = 21'b000000000000000100110;
		14'b10101000101100:	sigmoid = 21'b000000000000000100110;
		14'b10101000101101:	sigmoid = 21'b000000000000000100110;
		14'b10101000101110:	sigmoid = 21'b000000000000000100110;
		14'b10101000101111:	sigmoid = 21'b000000000000000100110;
		14'b10101000110000:	sigmoid = 21'b000000000000000100110;
		14'b10101000110001:	sigmoid = 21'b000000000000000100110;
		14'b10101000110010:	sigmoid = 21'b000000000000000100110;
		14'b10101000110011:	sigmoid = 21'b000000000000000100110;
		14'b10101000110100:	sigmoid = 21'b000000000000000100110;
		14'b10101000110101:	sigmoid = 21'b000000000000000100110;
		14'b10101000110110:	sigmoid = 21'b000000000000000100110;
		14'b10101000110111:	sigmoid = 21'b000000000000000100110;
		14'b10101000111000:	sigmoid = 21'b000000000000000100111;
		14'b10101000111001:	sigmoid = 21'b000000000000000100111;
		14'b10101000111010:	sigmoid = 21'b000000000000000100111;
		14'b10101000111011:	sigmoid = 21'b000000000000000100111;
		14'b10101000111100:	sigmoid = 21'b000000000000000100111;
		14'b10101000111101:	sigmoid = 21'b000000000000000100111;
		14'b10101000111110:	sigmoid = 21'b000000000000000100111;
		14'b10101000111111:	sigmoid = 21'b000000000000000100111;
		14'b10101001000000:	sigmoid = 21'b000000000000000100111;
		14'b10101001000001:	sigmoid = 21'b000000000000000100111;
		14'b10101001000010:	sigmoid = 21'b000000000000000100111;
		14'b10101001000011:	sigmoid = 21'b000000000000000100111;
		14'b10101001000100:	sigmoid = 21'b000000000000000101000;
		14'b10101001000101:	sigmoid = 21'b000000000000000101000;
		14'b10101001000110:	sigmoid = 21'b000000000000000101000;
		14'b10101001000111:	sigmoid = 21'b000000000000000101000;
		14'b10101001001000:	sigmoid = 21'b000000000000000101000;
		14'b10101001001001:	sigmoid = 21'b000000000000000101000;
		14'b10101001001010:	sigmoid = 21'b000000000000000101000;
		14'b10101001001011:	sigmoid = 21'b000000000000000101000;
		14'b10101001001100:	sigmoid = 21'b000000000000000101000;
		14'b10101001001101:	sigmoid = 21'b000000000000000101000;
		14'b10101001001110:	sigmoid = 21'b000000000000000101000;
		14'b10101001001111:	sigmoid = 21'b000000000000000101000;
		14'b10101001010000:	sigmoid = 21'b000000000000000101000;
		14'b10101001010001:	sigmoid = 21'b000000000000000101001;
		14'b10101001010010:	sigmoid = 21'b000000000000000101001;
		14'b10101001010011:	sigmoid = 21'b000000000000000101001;
		14'b10101001010100:	sigmoid = 21'b000000000000000101001;
		14'b10101001010101:	sigmoid = 21'b000000000000000101001;
		14'b10101001010110:	sigmoid = 21'b000000000000000101001;
		14'b10101001010111:	sigmoid = 21'b000000000000000101001;
		14'b10101001011000:	sigmoid = 21'b000000000000000101001;
		14'b10101001011001:	sigmoid = 21'b000000000000000101001;
		14'b10101001011010:	sigmoid = 21'b000000000000000101001;
		14'b10101001011011:	sigmoid = 21'b000000000000000101001;
		14'b10101001011100:	sigmoid = 21'b000000000000000101001;
		14'b10101001011101:	sigmoid = 21'b000000000000000101010;
		14'b10101001011110:	sigmoid = 21'b000000000000000101010;
		14'b10101001011111:	sigmoid = 21'b000000000000000101010;
		14'b10101001100000:	sigmoid = 21'b000000000000000101010;
		14'b10101001100001:	sigmoid = 21'b000000000000000101010;
		14'b10101001100010:	sigmoid = 21'b000000000000000101010;
		14'b10101001100011:	sigmoid = 21'b000000000000000101010;
		14'b10101001100100:	sigmoid = 21'b000000000000000101010;
		14'b10101001100101:	sigmoid = 21'b000000000000000101010;
		14'b10101001100110:	sigmoid = 21'b000000000000000101010;
		14'b10101001100111:	sigmoid = 21'b000000000000000101010;
		14'b10101001101000:	sigmoid = 21'b000000000000000101010;
		14'b10101001101001:	sigmoid = 21'b000000000000000101010;
		14'b10101001101010:	sigmoid = 21'b000000000000000101011;
		14'b10101001101011:	sigmoid = 21'b000000000000000101011;
		14'b10101001101100:	sigmoid = 21'b000000000000000101011;
		14'b10101001101101:	sigmoid = 21'b000000000000000101011;
		14'b10101001101110:	sigmoid = 21'b000000000000000101011;
		14'b10101001101111:	sigmoid = 21'b000000000000000101011;
		14'b10101001110000:	sigmoid = 21'b000000000000000101011;
		14'b10101001110001:	sigmoid = 21'b000000000000000101011;
		14'b10101001110010:	sigmoid = 21'b000000000000000101011;
		14'b10101001110011:	sigmoid = 21'b000000000000000101011;
		14'b10101001110100:	sigmoid = 21'b000000000000000101011;
		14'b10101001110101:	sigmoid = 21'b000000000000000101100;
		14'b10101001110110:	sigmoid = 21'b000000000000000101100;
		14'b10101001110111:	sigmoid = 21'b000000000000000101100;
		14'b10101001111000:	sigmoid = 21'b000000000000000101100;
		14'b10101001111001:	sigmoid = 21'b000000000000000101100;
		14'b10101001111010:	sigmoid = 21'b000000000000000101100;
		14'b10101001111011:	sigmoid = 21'b000000000000000101100;
		14'b10101001111100:	sigmoid = 21'b000000000000000101100;
		14'b10101001111101:	sigmoid = 21'b000000000000000101100;
		14'b10101001111110:	sigmoid = 21'b000000000000000101100;
		14'b10101001111111:	sigmoid = 21'b000000000000000101100;
		14'b10101010000000:	sigmoid = 21'b000000000000000101100;
		14'b10101010000001:	sigmoid = 21'b000000000000000101101;
		14'b10101010000010:	sigmoid = 21'b000000000000000101101;
		14'b10101010000011:	sigmoid = 21'b000000000000000101101;
		14'b10101010000100:	sigmoid = 21'b000000000000000101101;
		14'b10101010000101:	sigmoid = 21'b000000000000000101101;
		14'b10101010000110:	sigmoid = 21'b000000000000000101101;
		14'b10101010000111:	sigmoid = 21'b000000000000000101101;
		14'b10101010001000:	sigmoid = 21'b000000000000000101101;
		14'b10101010001001:	sigmoid = 21'b000000000000000101101;
		14'b10101010001010:	sigmoid = 21'b000000000000000101101;
		14'b10101010001011:	sigmoid = 21'b000000000000000101101;
		14'b10101010001100:	sigmoid = 21'b000000000000000101110;
		14'b10101010001101:	sigmoid = 21'b000000000000000101110;
		14'b10101010001110:	sigmoid = 21'b000000000000000101110;
		14'b10101010001111:	sigmoid = 21'b000000000000000101110;
		14'b10101010010000:	sigmoid = 21'b000000000000000101110;
		14'b10101010010001:	sigmoid = 21'b000000000000000101110;
		14'b10101010010010:	sigmoid = 21'b000000000000000101110;
		14'b10101010010011:	sigmoid = 21'b000000000000000101110;
		14'b10101010010100:	sigmoid = 21'b000000000000000101110;
		14'b10101010010101:	sigmoid = 21'b000000000000000101110;
		14'b10101010010110:	sigmoid = 21'b000000000000000101110;
		14'b10101010010111:	sigmoid = 21'b000000000000000101111;
		14'b10101010011000:	sigmoid = 21'b000000000000000101111;
		14'b10101010011001:	sigmoid = 21'b000000000000000101111;
		14'b10101010011010:	sigmoid = 21'b000000000000000101111;
		14'b10101010011011:	sigmoid = 21'b000000000000000101111;
		14'b10101010011100:	sigmoid = 21'b000000000000000101111;
		14'b10101010011101:	sigmoid = 21'b000000000000000101111;
		14'b10101010011110:	sigmoid = 21'b000000000000000101111;
		14'b10101010011111:	sigmoid = 21'b000000000000000101111;
		14'b10101010100000:	sigmoid = 21'b000000000000000101111;
		14'b10101010100001:	sigmoid = 21'b000000000000000101111;
		14'b10101010100010:	sigmoid = 21'b000000000000000110000;
		14'b10101010100011:	sigmoid = 21'b000000000000000110000;
		14'b10101010100100:	sigmoid = 21'b000000000000000110000;
		14'b10101010100101:	sigmoid = 21'b000000000000000110000;
		14'b10101010100110:	sigmoid = 21'b000000000000000110000;
		14'b10101010100111:	sigmoid = 21'b000000000000000110000;
		14'b10101010101000:	sigmoid = 21'b000000000000000110000;
		14'b10101010101001:	sigmoid = 21'b000000000000000110000;
		14'b10101010101010:	sigmoid = 21'b000000000000000110000;
		14'b10101010101011:	sigmoid = 21'b000000000000000110000;
		14'b10101010101100:	sigmoid = 21'b000000000000000110001;
		14'b10101010101101:	sigmoid = 21'b000000000000000110001;
		14'b10101010101110:	sigmoid = 21'b000000000000000110001;
		14'b10101010101111:	sigmoid = 21'b000000000000000110001;
		14'b10101010110000:	sigmoid = 21'b000000000000000110001;
		14'b10101010110001:	sigmoid = 21'b000000000000000110001;
		14'b10101010110010:	sigmoid = 21'b000000000000000110001;
		14'b10101010110011:	sigmoid = 21'b000000000000000110001;
		14'b10101010110100:	sigmoid = 21'b000000000000000110001;
		14'b10101010110101:	sigmoid = 21'b000000000000000110001;
		14'b10101010110110:	sigmoid = 21'b000000000000000110001;
		14'b10101010110111:	sigmoid = 21'b000000000000000110010;
		14'b10101010111000:	sigmoid = 21'b000000000000000110010;
		14'b10101010111001:	sigmoid = 21'b000000000000000110010;
		14'b10101010111010:	sigmoid = 21'b000000000000000110010;
		14'b10101010111011:	sigmoid = 21'b000000000000000110010;
		14'b10101010111100:	sigmoid = 21'b000000000000000110010;
		14'b10101010111101:	sigmoid = 21'b000000000000000110010;
		14'b10101010111110:	sigmoid = 21'b000000000000000110010;
		14'b10101010111111:	sigmoid = 21'b000000000000000110010;
		14'b10101011000000:	sigmoid = 21'b000000000000000110010;
		14'b10101011000001:	sigmoid = 21'b000000000000000110011;
		14'b10101011000010:	sigmoid = 21'b000000000000000110011;
		14'b10101011000011:	sigmoid = 21'b000000000000000110011;
		14'b10101011000100:	sigmoid = 21'b000000000000000110011;
		14'b10101011000101:	sigmoid = 21'b000000000000000110011;
		14'b10101011000110:	sigmoid = 21'b000000000000000110011;
		14'b10101011000111:	sigmoid = 21'b000000000000000110011;
		14'b10101011001000:	sigmoid = 21'b000000000000000110011;
		14'b10101011001001:	sigmoid = 21'b000000000000000110011;
		14'b10101011001010:	sigmoid = 21'b000000000000000110011;
		14'b10101011001011:	sigmoid = 21'b000000000000000110100;
		14'b10101011001100:	sigmoid = 21'b000000000000000110100;
		14'b10101011001101:	sigmoid = 21'b000000000000000110100;
		14'b10101011001110:	sigmoid = 21'b000000000000000110100;
		14'b10101011001111:	sigmoid = 21'b000000000000000110100;
		14'b10101011010000:	sigmoid = 21'b000000000000000110100;
		14'b10101011010001:	sigmoid = 21'b000000000000000110100;
		14'b10101011010010:	sigmoid = 21'b000000000000000110100;
		14'b10101011010011:	sigmoid = 21'b000000000000000110100;
		14'b10101011010100:	sigmoid = 21'b000000000000000110100;
		14'b10101011010101:	sigmoid = 21'b000000000000000110101;
		14'b10101011010110:	sigmoid = 21'b000000000000000110101;
		14'b10101011010111:	sigmoid = 21'b000000000000000110101;
		14'b10101011011000:	sigmoid = 21'b000000000000000110101;
		14'b10101011011001:	sigmoid = 21'b000000000000000110101;
		14'b10101011011010:	sigmoid = 21'b000000000000000110101;
		14'b10101011011011:	sigmoid = 21'b000000000000000110101;
		14'b10101011011100:	sigmoid = 21'b000000000000000110101;
		14'b10101011011101:	sigmoid = 21'b000000000000000110101;
		14'b10101011011110:	sigmoid = 21'b000000000000000110110;
		14'b10101011011111:	sigmoid = 21'b000000000000000110110;
		14'b10101011100000:	sigmoid = 21'b000000000000000110110;
		14'b10101011100001:	sigmoid = 21'b000000000000000110110;
		14'b10101011100010:	sigmoid = 21'b000000000000000110110;
		14'b10101011100011:	sigmoid = 21'b000000000000000110110;
		14'b10101011100100:	sigmoid = 21'b000000000000000110110;
		14'b10101011100101:	sigmoid = 21'b000000000000000110110;
		14'b10101011100110:	sigmoid = 21'b000000000000000110110;
		14'b10101011100111:	sigmoid = 21'b000000000000000110110;
		14'b10101011101000:	sigmoid = 21'b000000000000000110111;
		14'b10101011101001:	sigmoid = 21'b000000000000000110111;
		14'b10101011101010:	sigmoid = 21'b000000000000000110111;
		14'b10101011101011:	sigmoid = 21'b000000000000000110111;
		14'b10101011101100:	sigmoid = 21'b000000000000000110111;
		14'b10101011101101:	sigmoid = 21'b000000000000000110111;
		14'b10101011101110:	sigmoid = 21'b000000000000000110111;
		14'b10101011101111:	sigmoid = 21'b000000000000000110111;
		14'b10101011110000:	sigmoid = 21'b000000000000000110111;
		14'b10101011110001:	sigmoid = 21'b000000000000000111000;
		14'b10101011110010:	sigmoid = 21'b000000000000000111000;
		14'b10101011110011:	sigmoid = 21'b000000000000000111000;
		14'b10101011110100:	sigmoid = 21'b000000000000000111000;
		14'b10101011110101:	sigmoid = 21'b000000000000000111000;
		14'b10101011110110:	sigmoid = 21'b000000000000000111000;
		14'b10101011110111:	sigmoid = 21'b000000000000000111000;
		14'b10101011111000:	sigmoid = 21'b000000000000000111000;
		14'b10101011111001:	sigmoid = 21'b000000000000000111000;
		14'b10101011111010:	sigmoid = 21'b000000000000000111001;
		14'b10101011111011:	sigmoid = 21'b000000000000000111001;
		14'b10101011111100:	sigmoid = 21'b000000000000000111001;
		14'b10101011111101:	sigmoid = 21'b000000000000000111001;
		14'b10101011111110:	sigmoid = 21'b000000000000000111001;
		14'b10101011111111:	sigmoid = 21'b000000000000000111001;
		14'b10101100000000:	sigmoid = 21'b000000000000000111001;
		14'b10101100000001:	sigmoid = 21'b000000000000000111001;
		14'b10101100000010:	sigmoid = 21'b000000000000000111001;
		14'b10101100000011:	sigmoid = 21'b000000000000000111010;
		14'b10101100000100:	sigmoid = 21'b000000000000000111010;
		14'b10101100000101:	sigmoid = 21'b000000000000000111010;
		14'b10101100000110:	sigmoid = 21'b000000000000000111010;
		14'b10101100000111:	sigmoid = 21'b000000000000000111010;
		14'b10101100001000:	sigmoid = 21'b000000000000000111010;
		14'b10101100001001:	sigmoid = 21'b000000000000000111010;
		14'b10101100001010:	sigmoid = 21'b000000000000000111010;
		14'b10101100001011:	sigmoid = 21'b000000000000000111011;
		14'b10101100001100:	sigmoid = 21'b000000000000000111011;
		14'b10101100001101:	sigmoid = 21'b000000000000000111011;
		14'b10101100001110:	sigmoid = 21'b000000000000000111011;
		14'b10101100001111:	sigmoid = 21'b000000000000000111011;
		14'b10101100010000:	sigmoid = 21'b000000000000000111011;
		14'b10101100010001:	sigmoid = 21'b000000000000000111011;
		14'b10101100010010:	sigmoid = 21'b000000000000000111011;
		14'b10101100010011:	sigmoid = 21'b000000000000000111011;
		14'b10101100010100:	sigmoid = 21'b000000000000000111100;
		14'b10101100010101:	sigmoid = 21'b000000000000000111100;
		14'b10101100010110:	sigmoid = 21'b000000000000000111100;
		14'b10101100010111:	sigmoid = 21'b000000000000000111100;
		14'b10101100011000:	sigmoid = 21'b000000000000000111100;
		14'b10101100011001:	sigmoid = 21'b000000000000000111100;
		14'b10101100011010:	sigmoid = 21'b000000000000000111100;
		14'b10101100011011:	sigmoid = 21'b000000000000000111100;
		14'b10101100011100:	sigmoid = 21'b000000000000000111100;
		14'b10101100011101:	sigmoid = 21'b000000000000000111101;
		14'b10101100011110:	sigmoid = 21'b000000000000000111101;
		14'b10101100011111:	sigmoid = 21'b000000000000000111101;
		14'b10101100100000:	sigmoid = 21'b000000000000000111101;
		14'b10101100100001:	sigmoid = 21'b000000000000000111101;
		14'b10101100100010:	sigmoid = 21'b000000000000000111101;
		14'b10101100100011:	sigmoid = 21'b000000000000000111101;
		14'b10101100100100:	sigmoid = 21'b000000000000000111101;
		14'b10101100100101:	sigmoid = 21'b000000000000000111110;
		14'b10101100100110:	sigmoid = 21'b000000000000000111110;
		14'b10101100100111:	sigmoid = 21'b000000000000000111110;
		14'b10101100101000:	sigmoid = 21'b000000000000000111110;
		14'b10101100101001:	sigmoid = 21'b000000000000000111110;
		14'b10101100101010:	sigmoid = 21'b000000000000000111110;
		14'b10101100101011:	sigmoid = 21'b000000000000000111110;
		14'b10101100101100:	sigmoid = 21'b000000000000000111110;
		14'b10101100101101:	sigmoid = 21'b000000000000000111111;
		14'b10101100101110:	sigmoid = 21'b000000000000000111111;
		14'b10101100101111:	sigmoid = 21'b000000000000000111111;
		14'b10101100110000:	sigmoid = 21'b000000000000000111111;
		14'b10101100110001:	sigmoid = 21'b000000000000000111111;
		14'b10101100110010:	sigmoid = 21'b000000000000000111111;
		14'b10101100110011:	sigmoid = 21'b000000000000000111111;
		14'b10101100110100:	sigmoid = 21'b000000000000000111111;
		14'b10101100110101:	sigmoid = 21'b000000000000001000000;
		14'b10101100110110:	sigmoid = 21'b000000000000001000000;
		14'b10101100110111:	sigmoid = 21'b000000000000001000000;
		14'b10101100111000:	sigmoid = 21'b000000000000001000000;
		14'b10101100111001:	sigmoid = 21'b000000000000001000000;
		14'b10101100111010:	sigmoid = 21'b000000000000001000000;
		14'b10101100111011:	sigmoid = 21'b000000000000001000000;
		14'b10101100111100:	sigmoid = 21'b000000000000001000000;
		14'b10101100111101:	sigmoid = 21'b000000000000001000001;
		14'b10101100111110:	sigmoid = 21'b000000000000001000001;
		14'b10101100111111:	sigmoid = 21'b000000000000001000001;
		14'b10101101000000:	sigmoid = 21'b000000000000001000001;
		14'b10101101000001:	sigmoid = 21'b000000000000001000001;
		14'b10101101000010:	sigmoid = 21'b000000000000001000001;
		14'b10101101000011:	sigmoid = 21'b000000000000001000001;
		14'b10101101000100:	sigmoid = 21'b000000000000001000001;
		14'b10101101000101:	sigmoid = 21'b000000000000001000010;
		14'b10101101000110:	sigmoid = 21'b000000000000001000010;
		14'b10101101000111:	sigmoid = 21'b000000000000001000010;
		14'b10101101001000:	sigmoid = 21'b000000000000001000010;
		14'b10101101001001:	sigmoid = 21'b000000000000001000010;
		14'b10101101001010:	sigmoid = 21'b000000000000001000010;
		14'b10101101001011:	sigmoid = 21'b000000000000001000010;
		14'b10101101001100:	sigmoid = 21'b000000000000001000010;
		14'b10101101001101:	sigmoid = 21'b000000000000001000011;
		14'b10101101001110:	sigmoid = 21'b000000000000001000011;
		14'b10101101001111:	sigmoid = 21'b000000000000001000011;
		14'b10101101010000:	sigmoid = 21'b000000000000001000011;
		14'b10101101010001:	sigmoid = 21'b000000000000001000011;
		14'b10101101010010:	sigmoid = 21'b000000000000001000011;
		14'b10101101010011:	sigmoid = 21'b000000000000001000011;
		14'b10101101010100:	sigmoid = 21'b000000000000001000100;
		14'b10101101010101:	sigmoid = 21'b000000000000001000100;
		14'b10101101010110:	sigmoid = 21'b000000000000001000100;
		14'b10101101010111:	sigmoid = 21'b000000000000001000100;
		14'b10101101011000:	sigmoid = 21'b000000000000001000100;
		14'b10101101011001:	sigmoid = 21'b000000000000001000100;
		14'b10101101011010:	sigmoid = 21'b000000000000001000100;
		14'b10101101011011:	sigmoid = 21'b000000000000001000100;
		14'b10101101011100:	sigmoid = 21'b000000000000001000101;
		14'b10101101011101:	sigmoid = 21'b000000000000001000101;
		14'b10101101011110:	sigmoid = 21'b000000000000001000101;
		14'b10101101011111:	sigmoid = 21'b000000000000001000101;
		14'b10101101100000:	sigmoid = 21'b000000000000001000101;
		14'b10101101100001:	sigmoid = 21'b000000000000001000101;
		14'b10101101100010:	sigmoid = 21'b000000000000001000101;
		14'b10101101100011:	sigmoid = 21'b000000000000001000110;
		14'b10101101100100:	sigmoid = 21'b000000000000001000110;
		14'b10101101100101:	sigmoid = 21'b000000000000001000110;
		14'b10101101100110:	sigmoid = 21'b000000000000001000110;
		14'b10101101100111:	sigmoid = 21'b000000000000001000110;
		14'b10101101101000:	sigmoid = 21'b000000000000001000110;
		14'b10101101101001:	sigmoid = 21'b000000000000001000110;
		14'b10101101101010:	sigmoid = 21'b000000000000001000111;
		14'b10101101101011:	sigmoid = 21'b000000000000001000111;
		14'b10101101101100:	sigmoid = 21'b000000000000001000111;
		14'b10101101101101:	sigmoid = 21'b000000000000001000111;
		14'b10101101101110:	sigmoid = 21'b000000000000001000111;
		14'b10101101101111:	sigmoid = 21'b000000000000001000111;
		14'b10101101110000:	sigmoid = 21'b000000000000001000111;
		14'b10101101110001:	sigmoid = 21'b000000000000001001000;
		14'b10101101110010:	sigmoid = 21'b000000000000001001000;
		14'b10101101110011:	sigmoid = 21'b000000000000001001000;
		14'b10101101110100:	sigmoid = 21'b000000000000001001000;
		14'b10101101110101:	sigmoid = 21'b000000000000001001000;
		14'b10101101110110:	sigmoid = 21'b000000000000001001000;
		14'b10101101110111:	sigmoid = 21'b000000000000001001000;
		14'b10101101111000:	sigmoid = 21'b000000000000001001000;
		14'b10101101111001:	sigmoid = 21'b000000000000001001001;
		14'b10101101111010:	sigmoid = 21'b000000000000001001001;
		14'b10101101111011:	sigmoid = 21'b000000000000001001001;
		14'b10101101111100:	sigmoid = 21'b000000000000001001001;
		14'b10101101111101:	sigmoid = 21'b000000000000001001001;
		14'b10101101111110:	sigmoid = 21'b000000000000001001001;
		14'b10101101111111:	sigmoid = 21'b000000000000001001010;
		14'b10101110000000:	sigmoid = 21'b000000000000001001010;
		14'b10101110000001:	sigmoid = 21'b000000000000001001010;
		14'b10101110000010:	sigmoid = 21'b000000000000001001010;
		14'b10101110000011:	sigmoid = 21'b000000000000001001010;
		14'b10101110000100:	sigmoid = 21'b000000000000001001010;
		14'b10101110000101:	sigmoid = 21'b000000000000001001010;
		14'b10101110000110:	sigmoid = 21'b000000000000001001011;
		14'b10101110000111:	sigmoid = 21'b000000000000001001011;
		14'b10101110001000:	sigmoid = 21'b000000000000001001011;
		14'b10101110001001:	sigmoid = 21'b000000000000001001011;
		14'b10101110001010:	sigmoid = 21'b000000000000001001011;
		14'b10101110001011:	sigmoid = 21'b000000000000001001011;
		14'b10101110001100:	sigmoid = 21'b000000000000001001011;
		14'b10101110001101:	sigmoid = 21'b000000000000001001100;
		14'b10101110001110:	sigmoid = 21'b000000000000001001100;
		14'b10101110001111:	sigmoid = 21'b000000000000001001100;
		14'b10101110010000:	sigmoid = 21'b000000000000001001100;
		14'b10101110010001:	sigmoid = 21'b000000000000001001100;
		14'b10101110010010:	sigmoid = 21'b000000000000001001100;
		14'b10101110010011:	sigmoid = 21'b000000000000001001100;
		14'b10101110010100:	sigmoid = 21'b000000000000001001101;
		14'b10101110010101:	sigmoid = 21'b000000000000001001101;
		14'b10101110010110:	sigmoid = 21'b000000000000001001101;
		14'b10101110010111:	sigmoid = 21'b000000000000001001101;
		14'b10101110011000:	sigmoid = 21'b000000000000001001101;
		14'b10101110011001:	sigmoid = 21'b000000000000001001101;
		14'b10101110011010:	sigmoid = 21'b000000000000001001110;
		14'b10101110011011:	sigmoid = 21'b000000000000001001110;
		14'b10101110011100:	sigmoid = 21'b000000000000001001110;
		14'b10101110011101:	sigmoid = 21'b000000000000001001110;
		14'b10101110011110:	sigmoid = 21'b000000000000001001110;
		14'b10101110011111:	sigmoid = 21'b000000000000001001110;
		14'b10101110100000:	sigmoid = 21'b000000000000001001110;
		14'b10101110100001:	sigmoid = 21'b000000000000001001111;
		14'b10101110100010:	sigmoid = 21'b000000000000001001111;
		14'b10101110100011:	sigmoid = 21'b000000000000001001111;
		14'b10101110100100:	sigmoid = 21'b000000000000001001111;
		14'b10101110100101:	sigmoid = 21'b000000000000001001111;
		14'b10101110100110:	sigmoid = 21'b000000000000001001111;
		14'b10101110100111:	sigmoid = 21'b000000000000001010000;
		14'b10101110101000:	sigmoid = 21'b000000000000001010000;
		14'b10101110101001:	sigmoid = 21'b000000000000001010000;
		14'b10101110101010:	sigmoid = 21'b000000000000001010000;
		14'b10101110101011:	sigmoid = 21'b000000000000001010000;
		14'b10101110101100:	sigmoid = 21'b000000000000001010000;
		14'b10101110101101:	sigmoid = 21'b000000000000001010000;
		14'b10101110101110:	sigmoid = 21'b000000000000001010001;
		14'b10101110101111:	sigmoid = 21'b000000000000001010001;
		14'b10101110110000:	sigmoid = 21'b000000000000001010001;
		14'b10101110110001:	sigmoid = 21'b000000000000001010001;
		14'b10101110110010:	sigmoid = 21'b000000000000001010001;
		14'b10101110110011:	sigmoid = 21'b000000000000001010001;
		14'b10101110110100:	sigmoid = 21'b000000000000001010010;
		14'b10101110110101:	sigmoid = 21'b000000000000001010010;
		14'b10101110110110:	sigmoid = 21'b000000000000001010010;
		14'b10101110110111:	sigmoid = 21'b000000000000001010010;
		14'b10101110111000:	sigmoid = 21'b000000000000001010010;
		14'b10101110111001:	sigmoid = 21'b000000000000001010010;
		14'b10101110111010:	sigmoid = 21'b000000000000001010011;
		14'b10101110111011:	sigmoid = 21'b000000000000001010011;
		14'b10101110111100:	sigmoid = 21'b000000000000001010011;
		14'b10101110111101:	sigmoid = 21'b000000000000001010011;
		14'b10101110111110:	sigmoid = 21'b000000000000001010011;
		14'b10101110111111:	sigmoid = 21'b000000000000001010011;
		14'b10101111000000:	sigmoid = 21'b000000000000001010100;
		14'b10101111000001:	sigmoid = 21'b000000000000001010100;
		14'b10101111000010:	sigmoid = 21'b000000000000001010100;
		14'b10101111000011:	sigmoid = 21'b000000000000001010100;
		14'b10101111000100:	sigmoid = 21'b000000000000001010100;
		14'b10101111000101:	sigmoid = 21'b000000000000001010100;
		14'b10101111000110:	sigmoid = 21'b000000000000001010101;
		14'b10101111000111:	sigmoid = 21'b000000000000001010101;
		14'b10101111001000:	sigmoid = 21'b000000000000001010101;
		14'b10101111001001:	sigmoid = 21'b000000000000001010101;
		14'b10101111001010:	sigmoid = 21'b000000000000001010101;
		14'b10101111001011:	sigmoid = 21'b000000000000001010101;
		14'b10101111001100:	sigmoid = 21'b000000000000001010110;
		14'b10101111001101:	sigmoid = 21'b000000000000001010110;
		14'b10101111001110:	sigmoid = 21'b000000000000001010110;
		14'b10101111001111:	sigmoid = 21'b000000000000001010110;
		14'b10101111010000:	sigmoid = 21'b000000000000001010110;
		14'b10101111010001:	sigmoid = 21'b000000000000001010110;
		14'b10101111010010:	sigmoid = 21'b000000000000001010111;
		14'b10101111010011:	sigmoid = 21'b000000000000001010111;
		14'b10101111010100:	sigmoid = 21'b000000000000001010111;
		14'b10101111010101:	sigmoid = 21'b000000000000001010111;
		14'b10101111010110:	sigmoid = 21'b000000000000001010111;
		14'b10101111010111:	sigmoid = 21'b000000000000001010111;
		14'b10101111011000:	sigmoid = 21'b000000000000001011000;
		14'b10101111011001:	sigmoid = 21'b000000000000001011000;
		14'b10101111011010:	sigmoid = 21'b000000000000001011000;
		14'b10101111011011:	sigmoid = 21'b000000000000001011000;
		14'b10101111011100:	sigmoid = 21'b000000000000001011000;
		14'b10101111011101:	sigmoid = 21'b000000000000001011000;
		14'b10101111011110:	sigmoid = 21'b000000000000001011001;
		14'b10101111011111:	sigmoid = 21'b000000000000001011001;
		14'b10101111100000:	sigmoid = 21'b000000000000001011001;
		14'b10101111100001:	sigmoid = 21'b000000000000001011001;
		14'b10101111100010:	sigmoid = 21'b000000000000001011001;
		14'b10101111100011:	sigmoid = 21'b000000000000001011001;
		14'b10101111100100:	sigmoid = 21'b000000000000001011010;
		14'b10101111100101:	sigmoid = 21'b000000000000001011010;
		14'b10101111100110:	sigmoid = 21'b000000000000001011010;
		14'b10101111100111:	sigmoid = 21'b000000000000001011010;
		14'b10101111101000:	sigmoid = 21'b000000000000001011010;
		14'b10101111101001:	sigmoid = 21'b000000000000001011011;
		14'b10101111101010:	sigmoid = 21'b000000000000001011011;
		14'b10101111101011:	sigmoid = 21'b000000000000001011011;
		14'b10101111101100:	sigmoid = 21'b000000000000001011011;
		14'b10101111101101:	sigmoid = 21'b000000000000001011011;
		14'b10101111101110:	sigmoid = 21'b000000000000001011011;
		14'b10101111101111:	sigmoid = 21'b000000000000001011100;
		14'b10101111110000:	sigmoid = 21'b000000000000001011100;
		14'b10101111110001:	sigmoid = 21'b000000000000001011100;
		14'b10101111110010:	sigmoid = 21'b000000000000001011100;
		14'b10101111110011:	sigmoid = 21'b000000000000001011100;
		14'b10101111110100:	sigmoid = 21'b000000000000001011101;
		14'b10101111110101:	sigmoid = 21'b000000000000001011101;
		14'b10101111110110:	sigmoid = 21'b000000000000001011101;
		14'b10101111110111:	sigmoid = 21'b000000000000001011101;
		14'b10101111111000:	sigmoid = 21'b000000000000001011101;
		14'b10101111111001:	sigmoid = 21'b000000000000001011101;
		14'b10101111111010:	sigmoid = 21'b000000000000001011110;
		14'b10101111111011:	sigmoid = 21'b000000000000001011110;
		14'b10101111111100:	sigmoid = 21'b000000000000001011110;
		14'b10101111111101:	sigmoid = 21'b000000000000001011110;
		14'b10101111111110:	sigmoid = 21'b000000000000001011110;
		14'b10101111111111:	sigmoid = 21'b000000000000001011111;
		14'b10110000000000:	sigmoid = 21'b000000000000001011111;
		14'b10110000000001:	sigmoid = 21'b000000000000001011111;
		14'b10110000000010:	sigmoid = 21'b000000000000001011111;
		14'b10110000000011:	sigmoid = 21'b000000000000001011111;
		14'b10110000000100:	sigmoid = 21'b000000000000001011111;
		14'b10110000000101:	sigmoid = 21'b000000000000001100000;
		14'b10110000000110:	sigmoid = 21'b000000000000001100000;
		14'b10110000000111:	sigmoid = 21'b000000000000001100000;
		14'b10110000001000:	sigmoid = 21'b000000000000001100000;
		14'b10110000001001:	sigmoid = 21'b000000000000001100000;
		14'b10110000001010:	sigmoid = 21'b000000000000001100001;
		14'b10110000001011:	sigmoid = 21'b000000000000001100001;
		14'b10110000001100:	sigmoid = 21'b000000000000001100001;
		14'b10110000001101:	sigmoid = 21'b000000000000001100001;
		14'b10110000001110:	sigmoid = 21'b000000000000001100001;
		14'b10110000001111:	sigmoid = 21'b000000000000001100010;
		14'b10110000010000:	sigmoid = 21'b000000000000001100010;
		14'b10110000010001:	sigmoid = 21'b000000000000001100010;
		14'b10110000010010:	sigmoid = 21'b000000000000001100010;
		14'b10110000010011:	sigmoid = 21'b000000000000001100010;
		14'b10110000010100:	sigmoid = 21'b000000000000001100010;
		14'b10110000010101:	sigmoid = 21'b000000000000001100011;
		14'b10110000010110:	sigmoid = 21'b000000000000001100011;
		14'b10110000010111:	sigmoid = 21'b000000000000001100011;
		14'b10110000011000:	sigmoid = 21'b000000000000001100011;
		14'b10110000011001:	sigmoid = 21'b000000000000001100011;
		14'b10110000011010:	sigmoid = 21'b000000000000001100100;
		14'b10110000011011:	sigmoid = 21'b000000000000001100100;
		14'b10110000011100:	sigmoid = 21'b000000000000001100100;
		14'b10110000011101:	sigmoid = 21'b000000000000001100100;
		14'b10110000011110:	sigmoid = 21'b000000000000001100100;
		14'b10110000011111:	sigmoid = 21'b000000000000001100101;
		14'b10110000100000:	sigmoid = 21'b000000000000001100101;
		14'b10110000100001:	sigmoid = 21'b000000000000001100101;
		14'b10110000100010:	sigmoid = 21'b000000000000001100101;
		14'b10110000100011:	sigmoid = 21'b000000000000001100101;
		14'b10110000100100:	sigmoid = 21'b000000000000001100110;
		14'b10110000100101:	sigmoid = 21'b000000000000001100110;
		14'b10110000100110:	sigmoid = 21'b000000000000001100110;
		14'b10110000100111:	sigmoid = 21'b000000000000001100110;
		14'b10110000101000:	sigmoid = 21'b000000000000001100110;
		14'b10110000101001:	sigmoid = 21'b000000000000001100111;
		14'b10110000101010:	sigmoid = 21'b000000000000001100111;
		14'b10110000101011:	sigmoid = 21'b000000000000001100111;
		14'b10110000101100:	sigmoid = 21'b000000000000001100111;
		14'b10110000101101:	sigmoid = 21'b000000000000001100111;
		14'b10110000101110:	sigmoid = 21'b000000000000001101000;
		14'b10110000101111:	sigmoid = 21'b000000000000001101000;
		14'b10110000110000:	sigmoid = 21'b000000000000001101000;
		14'b10110000110001:	sigmoid = 21'b000000000000001101000;
		14'b10110000110010:	sigmoid = 21'b000000000000001101000;
		14'b10110000110011:	sigmoid = 21'b000000000000001101001;
		14'b10110000110100:	sigmoid = 21'b000000000000001101001;
		14'b10110000110101:	sigmoid = 21'b000000000000001101001;
		14'b10110000110110:	sigmoid = 21'b000000000000001101001;
		14'b10110000110111:	sigmoid = 21'b000000000000001101010;
		14'b10110000111000:	sigmoid = 21'b000000000000001101010;
		14'b10110000111001:	sigmoid = 21'b000000000000001101010;
		14'b10110000111010:	sigmoid = 21'b000000000000001101010;
		14'b10110000111011:	sigmoid = 21'b000000000000001101010;
		14'b10110000111100:	sigmoid = 21'b000000000000001101011;
		14'b10110000111101:	sigmoid = 21'b000000000000001101011;
		14'b10110000111110:	sigmoid = 21'b000000000000001101011;
		14'b10110000111111:	sigmoid = 21'b000000000000001101011;
		14'b10110001000000:	sigmoid = 21'b000000000000001101011;
		14'b10110001000001:	sigmoid = 21'b000000000000001101100;
		14'b10110001000010:	sigmoid = 21'b000000000000001101100;
		14'b10110001000011:	sigmoid = 21'b000000000000001101100;
		14'b10110001000100:	sigmoid = 21'b000000000000001101100;
		14'b10110001000101:	sigmoid = 21'b000000000000001101100;
		14'b10110001000110:	sigmoid = 21'b000000000000001101101;
		14'b10110001000111:	sigmoid = 21'b000000000000001101101;
		14'b10110001001000:	sigmoid = 21'b000000000000001101101;
		14'b10110001001001:	sigmoid = 21'b000000000000001101101;
		14'b10110001001010:	sigmoid = 21'b000000000000001101110;
		14'b10110001001011:	sigmoid = 21'b000000000000001101110;
		14'b10110001001100:	sigmoid = 21'b000000000000001101110;
		14'b10110001001101:	sigmoid = 21'b000000000000001101110;
		14'b10110001001110:	sigmoid = 21'b000000000000001101110;
		14'b10110001001111:	sigmoid = 21'b000000000000001101111;
		14'b10110001010000:	sigmoid = 21'b000000000000001101111;
		14'b10110001010001:	sigmoid = 21'b000000000000001101111;
		14'b10110001010010:	sigmoid = 21'b000000000000001101111;
		14'b10110001010011:	sigmoid = 21'b000000000000001101111;
		14'b10110001010100:	sigmoid = 21'b000000000000001110000;
		14'b10110001010101:	sigmoid = 21'b000000000000001110000;
		14'b10110001010110:	sigmoid = 21'b000000000000001110000;
		14'b10110001010111:	sigmoid = 21'b000000000000001110000;
		14'b10110001011000:	sigmoid = 21'b000000000000001110001;
		14'b10110001011001:	sigmoid = 21'b000000000000001110001;
		14'b10110001011010:	sigmoid = 21'b000000000000001110001;
		14'b10110001011011:	sigmoid = 21'b000000000000001110001;
		14'b10110001011100:	sigmoid = 21'b000000000000001110001;
		14'b10110001011101:	sigmoid = 21'b000000000000001110010;
		14'b10110001011110:	sigmoid = 21'b000000000000001110010;
		14'b10110001011111:	sigmoid = 21'b000000000000001110010;
		14'b10110001100000:	sigmoid = 21'b000000000000001110010;
		14'b10110001100001:	sigmoid = 21'b000000000000001110011;
		14'b10110001100010:	sigmoid = 21'b000000000000001110011;
		14'b10110001100011:	sigmoid = 21'b000000000000001110011;
		14'b10110001100100:	sigmoid = 21'b000000000000001110011;
		14'b10110001100101:	sigmoid = 21'b000000000000001110011;
		14'b10110001100110:	sigmoid = 21'b000000000000001110100;
		14'b10110001100111:	sigmoid = 21'b000000000000001110100;
		14'b10110001101000:	sigmoid = 21'b000000000000001110100;
		14'b10110001101001:	sigmoid = 21'b000000000000001110100;
		14'b10110001101010:	sigmoid = 21'b000000000000001110101;
		14'b10110001101011:	sigmoid = 21'b000000000000001110101;
		14'b10110001101100:	sigmoid = 21'b000000000000001110101;
		14'b10110001101101:	sigmoid = 21'b000000000000001110101;
		14'b10110001101110:	sigmoid = 21'b000000000000001110110;
		14'b10110001101111:	sigmoid = 21'b000000000000001110110;
		14'b10110001110000:	sigmoid = 21'b000000000000001110110;
		14'b10110001110001:	sigmoid = 21'b000000000000001110110;
		14'b10110001110010:	sigmoid = 21'b000000000000001110110;
		14'b10110001110011:	sigmoid = 21'b000000000000001110111;
		14'b10110001110100:	sigmoid = 21'b000000000000001110111;
		14'b10110001110101:	sigmoid = 21'b000000000000001110111;
		14'b10110001110110:	sigmoid = 21'b000000000000001110111;
		14'b10110001110111:	sigmoid = 21'b000000000000001111000;
		14'b10110001111000:	sigmoid = 21'b000000000000001111000;
		14'b10110001111001:	sigmoid = 21'b000000000000001111000;
		14'b10110001111010:	sigmoid = 21'b000000000000001111000;
		14'b10110001111011:	sigmoid = 21'b000000000000001111001;
		14'b10110001111100:	sigmoid = 21'b000000000000001111001;
		14'b10110001111101:	sigmoid = 21'b000000000000001111001;
		14'b10110001111110:	sigmoid = 21'b000000000000001111001;
		14'b10110001111111:	sigmoid = 21'b000000000000001111010;
		14'b10110010000000:	sigmoid = 21'b000000000000001111010;
		14'b10110010000001:	sigmoid = 21'b000000000000001111010;
		14'b10110010000010:	sigmoid = 21'b000000000000001111010;
		14'b10110010000011:	sigmoid = 21'b000000000000001111010;
		14'b10110010000100:	sigmoid = 21'b000000000000001111011;
		14'b10110010000101:	sigmoid = 21'b000000000000001111011;
		14'b10110010000110:	sigmoid = 21'b000000000000001111011;
		14'b10110010000111:	sigmoid = 21'b000000000000001111011;
		14'b10110010001000:	sigmoid = 21'b000000000000001111100;
		14'b10110010001001:	sigmoid = 21'b000000000000001111100;
		14'b10110010001010:	sigmoid = 21'b000000000000001111100;
		14'b10110010001011:	sigmoid = 21'b000000000000001111100;
		14'b10110010001100:	sigmoid = 21'b000000000000001111101;
		14'b10110010001101:	sigmoid = 21'b000000000000001111101;
		14'b10110010001110:	sigmoid = 21'b000000000000001111101;
		14'b10110010001111:	sigmoid = 21'b000000000000001111101;
		14'b10110010010000:	sigmoid = 21'b000000000000001111110;
		14'b10110010010001:	sigmoid = 21'b000000000000001111110;
		14'b10110010010010:	sigmoid = 21'b000000000000001111110;
		14'b10110010010011:	sigmoid = 21'b000000000000001111110;
		14'b10110010010100:	sigmoid = 21'b000000000000001111111;
		14'b10110010010101:	sigmoid = 21'b000000000000001111111;
		14'b10110010010110:	sigmoid = 21'b000000000000001111111;
		14'b10110010010111:	sigmoid = 21'b000000000000001111111;
		14'b10110010011000:	sigmoid = 21'b000000000000010000000;
		14'b10110010011001:	sigmoid = 21'b000000000000010000000;
		14'b10110010011010:	sigmoid = 21'b000000000000010000000;
		14'b10110010011011:	sigmoid = 21'b000000000000010000000;
		14'b10110010011100:	sigmoid = 21'b000000000000010000001;
		14'b10110010011101:	sigmoid = 21'b000000000000010000001;
		14'b10110010011110:	sigmoid = 21'b000000000000010000001;
		14'b10110010011111:	sigmoid = 21'b000000000000010000001;
		14'b10110010100000:	sigmoid = 21'b000000000000010000010;
		14'b10110010100001:	sigmoid = 21'b000000000000010000010;
		14'b10110010100010:	sigmoid = 21'b000000000000010000010;
		14'b10110010100011:	sigmoid = 21'b000000000000010000010;
		14'b10110010100100:	sigmoid = 21'b000000000000010000011;
		14'b10110010100101:	sigmoid = 21'b000000000000010000011;
		14'b10110010100110:	sigmoid = 21'b000000000000010000011;
		14'b10110010100111:	sigmoid = 21'b000000000000010000011;
		14'b10110010101000:	sigmoid = 21'b000000000000010000100;
		14'b10110010101001:	sigmoid = 21'b000000000000010000100;
		14'b10110010101010:	sigmoid = 21'b000000000000010000100;
		14'b10110010101011:	sigmoid = 21'b000000000000010000100;
		14'b10110010101100:	sigmoid = 21'b000000000000010000101;
		14'b10110010101101:	sigmoid = 21'b000000000000010000101;
		14'b10110010101110:	sigmoid = 21'b000000000000010000101;
		14'b10110010101111:	sigmoid = 21'b000000000000010000101;
		14'b10110010110000:	sigmoid = 21'b000000000000010000110;
		14'b10110010110001:	sigmoid = 21'b000000000000010000110;
		14'b10110010110010:	sigmoid = 21'b000000000000010000110;
		14'b10110010110011:	sigmoid = 21'b000000000000010000111;
		14'b10110010110100:	sigmoid = 21'b000000000000010000111;
		14'b10110010110101:	sigmoid = 21'b000000000000010000111;
		14'b10110010110110:	sigmoid = 21'b000000000000010000111;
		14'b10110010110111:	sigmoid = 21'b000000000000010001000;
		14'b10110010111000:	sigmoid = 21'b000000000000010001000;
		14'b10110010111001:	sigmoid = 21'b000000000000010001000;
		14'b10110010111010:	sigmoid = 21'b000000000000010001000;
		14'b10110010111011:	sigmoid = 21'b000000000000010001001;
		14'b10110010111100:	sigmoid = 21'b000000000000010001001;
		14'b10110010111101:	sigmoid = 21'b000000000000010001001;
		14'b10110010111110:	sigmoid = 21'b000000000000010001001;
		14'b10110010111111:	sigmoid = 21'b000000000000010001010;
		14'b10110011000000:	sigmoid = 21'b000000000000010001010;
		14'b10110011000001:	sigmoid = 21'b000000000000010001010;
		14'b10110011000010:	sigmoid = 21'b000000000000010001011;
		14'b10110011000011:	sigmoid = 21'b000000000000010001011;
		14'b10110011000100:	sigmoid = 21'b000000000000010001011;
		14'b10110011000101:	sigmoid = 21'b000000000000010001011;
		14'b10110011000110:	sigmoid = 21'b000000000000010001100;
		14'b10110011000111:	sigmoid = 21'b000000000000010001100;
		14'b10110011001000:	sigmoid = 21'b000000000000010001100;
		14'b10110011001001:	sigmoid = 21'b000000000000010001100;
		14'b10110011001010:	sigmoid = 21'b000000000000010001101;
		14'b10110011001011:	sigmoid = 21'b000000000000010001101;
		14'b10110011001100:	sigmoid = 21'b000000000000010001101;
		14'b10110011001101:	sigmoid = 21'b000000000000010001110;
		14'b10110011001110:	sigmoid = 21'b000000000000010001110;
		14'b10110011001111:	sigmoid = 21'b000000000000010001110;
		14'b10110011010000:	sigmoid = 21'b000000000000010001110;
		14'b10110011010001:	sigmoid = 21'b000000000000010001111;
		14'b10110011010010:	sigmoid = 21'b000000000000010001111;
		14'b10110011010011:	sigmoid = 21'b000000000000010001111;
		14'b10110011010100:	sigmoid = 21'b000000000000010010000;
		14'b10110011010101:	sigmoid = 21'b000000000000010010000;
		14'b10110011010110:	sigmoid = 21'b000000000000010010000;
		14'b10110011010111:	sigmoid = 21'b000000000000010010000;
		14'b10110011011000:	sigmoid = 21'b000000000000010010001;
		14'b10110011011001:	sigmoid = 21'b000000000000010010001;
		14'b10110011011010:	sigmoid = 21'b000000000000010010001;
		14'b10110011011011:	sigmoid = 21'b000000000000010010010;
		14'b10110011011100:	sigmoid = 21'b000000000000010010010;
		14'b10110011011101:	sigmoid = 21'b000000000000010010010;
		14'b10110011011110:	sigmoid = 21'b000000000000010010010;
		14'b10110011011111:	sigmoid = 21'b000000000000010010011;
		14'b10110011100000:	sigmoid = 21'b000000000000010010011;
		14'b10110011100001:	sigmoid = 21'b000000000000010010011;
		14'b10110011100010:	sigmoid = 21'b000000000000010010100;
		14'b10110011100011:	sigmoid = 21'b000000000000010010100;
		14'b10110011100100:	sigmoid = 21'b000000000000010010100;
		14'b10110011100101:	sigmoid = 21'b000000000000010010100;
		14'b10110011100110:	sigmoid = 21'b000000000000010010101;
		14'b10110011100111:	sigmoid = 21'b000000000000010010101;
		14'b10110011101000:	sigmoid = 21'b000000000000010010101;
		14'b10110011101001:	sigmoid = 21'b000000000000010010110;
		14'b10110011101010:	sigmoid = 21'b000000000000010010110;
		14'b10110011101011:	sigmoid = 21'b000000000000010010110;
		14'b10110011101100:	sigmoid = 21'b000000000000010010110;
		14'b10110011101101:	sigmoid = 21'b000000000000010010111;
		14'b10110011101110:	sigmoid = 21'b000000000000010010111;
		14'b10110011101111:	sigmoid = 21'b000000000000010010111;
		14'b10110011110000:	sigmoid = 21'b000000000000010011000;
		14'b10110011110001:	sigmoid = 21'b000000000000010011000;
		14'b10110011110010:	sigmoid = 21'b000000000000010011000;
		14'b10110011110011:	sigmoid = 21'b000000000000010011001;
		14'b10110011110100:	sigmoid = 21'b000000000000010011001;
		14'b10110011110101:	sigmoid = 21'b000000000000010011001;
		14'b10110011110110:	sigmoid = 21'b000000000000010011001;
		14'b10110011110111:	sigmoid = 21'b000000000000010011010;
		14'b10110011111000:	sigmoid = 21'b000000000000010011010;
		14'b10110011111001:	sigmoid = 21'b000000000000010011010;
		14'b10110011111010:	sigmoid = 21'b000000000000010011011;
		14'b10110011111011:	sigmoid = 21'b000000000000010011011;
		14'b10110011111100:	sigmoid = 21'b000000000000010011011;
		14'b10110011111101:	sigmoid = 21'b000000000000010011100;
		14'b10110011111110:	sigmoid = 21'b000000000000010011100;
		14'b10110011111111:	sigmoid = 21'b000000000000010011100;
		14'b10110100000000:	sigmoid = 21'b000000000000010011100;
		14'b10110100000001:	sigmoid = 21'b000000000000010011101;
		14'b10110100000010:	sigmoid = 21'b000000000000010011101;
		14'b10110100000011:	sigmoid = 21'b000000000000010011101;
		14'b10110100000100:	sigmoid = 21'b000000000000010011110;
		14'b10110100000101:	sigmoid = 21'b000000000000010011110;
		14'b10110100000110:	sigmoid = 21'b000000000000010011110;
		14'b10110100000111:	sigmoid = 21'b000000000000010011111;
		14'b10110100001000:	sigmoid = 21'b000000000000010011111;
		14'b10110100001001:	sigmoid = 21'b000000000000010011111;
		14'b10110100001010:	sigmoid = 21'b000000000000010100000;
		14'b10110100001011:	sigmoid = 21'b000000000000010100000;
		14'b10110100001100:	sigmoid = 21'b000000000000010100000;
		14'b10110100001101:	sigmoid = 21'b000000000000010100001;
		14'b10110100001110:	sigmoid = 21'b000000000000010100001;
		14'b10110100001111:	sigmoid = 21'b000000000000010100001;
		14'b10110100010000:	sigmoid = 21'b000000000000010100001;
		14'b10110100010001:	sigmoid = 21'b000000000000010100010;
		14'b10110100010010:	sigmoid = 21'b000000000000010100010;
		14'b10110100010011:	sigmoid = 21'b000000000000010100010;
		14'b10110100010100:	sigmoid = 21'b000000000000010100011;
		14'b10110100010101:	sigmoid = 21'b000000000000010100011;
		14'b10110100010110:	sigmoid = 21'b000000000000010100011;
		14'b10110100010111:	sigmoid = 21'b000000000000010100100;
		14'b10110100011000:	sigmoid = 21'b000000000000010100100;
		14'b10110100011001:	sigmoid = 21'b000000000000010100100;
		14'b10110100011010:	sigmoid = 21'b000000000000010100101;
		14'b10110100011011:	sigmoid = 21'b000000000000010100101;
		14'b10110100011100:	sigmoid = 21'b000000000000010100101;
		14'b10110100011101:	sigmoid = 21'b000000000000010100110;
		14'b10110100011110:	sigmoid = 21'b000000000000010100110;
		14'b10110100011111:	sigmoid = 21'b000000000000010100110;
		14'b10110100100000:	sigmoid = 21'b000000000000010100111;
		14'b10110100100001:	sigmoid = 21'b000000000000010100111;
		14'b10110100100010:	sigmoid = 21'b000000000000010100111;
		14'b10110100100011:	sigmoid = 21'b000000000000010101000;
		14'b10110100100100:	sigmoid = 21'b000000000000010101000;
		14'b10110100100101:	sigmoid = 21'b000000000000010101000;
		14'b10110100100110:	sigmoid = 21'b000000000000010101001;
		14'b10110100100111:	sigmoid = 21'b000000000000010101001;
		14'b10110100101000:	sigmoid = 21'b000000000000010101001;
		14'b10110100101001:	sigmoid = 21'b000000000000010101010;
		14'b10110100101010:	sigmoid = 21'b000000000000010101010;
		14'b10110100101011:	sigmoid = 21'b000000000000010101010;
		14'b10110100101100:	sigmoid = 21'b000000000000010101011;
		14'b10110100101101:	sigmoid = 21'b000000000000010101011;
		14'b10110100101110:	sigmoid = 21'b000000000000010101011;
		14'b10110100101111:	sigmoid = 21'b000000000000010101100;
		14'b10110100110000:	sigmoid = 21'b000000000000010101100;
		14'b10110100110001:	sigmoid = 21'b000000000000010101100;
		14'b10110100110010:	sigmoid = 21'b000000000000010101101;
		14'b10110100110011:	sigmoid = 21'b000000000000010101101;
		14'b10110100110100:	sigmoid = 21'b000000000000010101101;
		14'b10110100110101:	sigmoid = 21'b000000000000010101110;
		14'b10110100110110:	sigmoid = 21'b000000000000010101110;
		14'b10110100110111:	sigmoid = 21'b000000000000010101110;
		14'b10110100111000:	sigmoid = 21'b000000000000010101111;
		14'b10110100111001:	sigmoid = 21'b000000000000010101111;
		14'b10110100111010:	sigmoid = 21'b000000000000010101111;
		14'b10110100111011:	sigmoid = 21'b000000000000010110000;
		14'b10110100111100:	sigmoid = 21'b000000000000010110000;
		14'b10110100111101:	sigmoid = 21'b000000000000010110000;
		14'b10110100111110:	sigmoid = 21'b000000000000010110001;
		14'b10110100111111:	sigmoid = 21'b000000000000010110001;
		14'b10110101000000:	sigmoid = 21'b000000000000010110001;
		14'b10110101000001:	sigmoid = 21'b000000000000010110010;
		14'b10110101000010:	sigmoid = 21'b000000000000010110010;
		14'b10110101000011:	sigmoid = 21'b000000000000010110010;
		14'b10110101000100:	sigmoid = 21'b000000000000010110011;
		14'b10110101000101:	sigmoid = 21'b000000000000010110011;
		14'b10110101000110:	sigmoid = 21'b000000000000010110011;
		14'b10110101000111:	sigmoid = 21'b000000000000010110100;
		14'b10110101001000:	sigmoid = 21'b000000000000010110100;
		14'b10110101001001:	sigmoid = 21'b000000000000010110101;
		14'b10110101001010:	sigmoid = 21'b000000000000010110101;
		14'b10110101001011:	sigmoid = 21'b000000000000010110101;
		14'b10110101001100:	sigmoid = 21'b000000000000010110110;
		14'b10110101001101:	sigmoid = 21'b000000000000010110110;
		14'b10110101001110:	sigmoid = 21'b000000000000010110110;
		14'b10110101001111:	sigmoid = 21'b000000000000010110111;
		14'b10110101010000:	sigmoid = 21'b000000000000010110111;
		14'b10110101010001:	sigmoid = 21'b000000000000010110111;
		14'b10110101010010:	sigmoid = 21'b000000000000010111000;
		14'b10110101010011:	sigmoid = 21'b000000000000010111000;
		14'b10110101010100:	sigmoid = 21'b000000000000010111000;
		14'b10110101010101:	sigmoid = 21'b000000000000010111001;
		14'b10110101010110:	sigmoid = 21'b000000000000010111001;
		14'b10110101010111:	sigmoid = 21'b000000000000010111010;
		14'b10110101011000:	sigmoid = 21'b000000000000010111010;
		14'b10110101011001:	sigmoid = 21'b000000000000010111010;
		14'b10110101011010:	sigmoid = 21'b000000000000010111011;
		14'b10110101011011:	sigmoid = 21'b000000000000010111011;
		14'b10110101011100:	sigmoid = 21'b000000000000010111011;
		14'b10110101011101:	sigmoid = 21'b000000000000010111100;
		14'b10110101011110:	sigmoid = 21'b000000000000010111100;
		14'b10110101011111:	sigmoid = 21'b000000000000010111100;
		14'b10110101100000:	sigmoid = 21'b000000000000010111101;
		14'b10110101100001:	sigmoid = 21'b000000000000010111101;
		14'b10110101100010:	sigmoid = 21'b000000000000010111110;
		14'b10110101100011:	sigmoid = 21'b000000000000010111110;
		14'b10110101100100:	sigmoid = 21'b000000000000010111110;
		14'b10110101100101:	sigmoid = 21'b000000000000010111111;
		14'b10110101100110:	sigmoid = 21'b000000000000010111111;
		14'b10110101100111:	sigmoid = 21'b000000000000010111111;
		14'b10110101101000:	sigmoid = 21'b000000000000011000000;
		14'b10110101101001:	sigmoid = 21'b000000000000011000000;
		14'b10110101101010:	sigmoid = 21'b000000000000011000001;
		14'b10110101101011:	sigmoid = 21'b000000000000011000001;
		14'b10110101101100:	sigmoid = 21'b000000000000011000001;
		14'b10110101101101:	sigmoid = 21'b000000000000011000010;
		14'b10110101101110:	sigmoid = 21'b000000000000011000010;
		14'b10110101101111:	sigmoid = 21'b000000000000011000010;
		14'b10110101110000:	sigmoid = 21'b000000000000011000011;
		14'b10110101110001:	sigmoid = 21'b000000000000011000011;
		14'b10110101110010:	sigmoid = 21'b000000000000011000100;
		14'b10110101110011:	sigmoid = 21'b000000000000011000100;
		14'b10110101110100:	sigmoid = 21'b000000000000011000100;
		14'b10110101110101:	sigmoid = 21'b000000000000011000101;
		14'b10110101110110:	sigmoid = 21'b000000000000011000101;
		14'b10110101110111:	sigmoid = 21'b000000000000011000110;
		14'b10110101111000:	sigmoid = 21'b000000000000011000110;
		14'b10110101111001:	sigmoid = 21'b000000000000011000110;
		14'b10110101111010:	sigmoid = 21'b000000000000011000111;
		14'b10110101111011:	sigmoid = 21'b000000000000011000111;
		14'b10110101111100:	sigmoid = 21'b000000000000011000111;
		14'b10110101111101:	sigmoid = 21'b000000000000011001000;
		14'b10110101111110:	sigmoid = 21'b000000000000011001000;
		14'b10110101111111:	sigmoid = 21'b000000000000011001001;
		14'b10110110000000:	sigmoid = 21'b000000000000011001001;
		14'b10110110000001:	sigmoid = 21'b000000000000011001001;
		14'b10110110000010:	sigmoid = 21'b000000000000011001010;
		14'b10110110000011:	sigmoid = 21'b000000000000011001010;
		14'b10110110000100:	sigmoid = 21'b000000000000011001011;
		14'b10110110000101:	sigmoid = 21'b000000000000011001011;
		14'b10110110000110:	sigmoid = 21'b000000000000011001011;
		14'b10110110000111:	sigmoid = 21'b000000000000011001100;
		14'b10110110001000:	sigmoid = 21'b000000000000011001100;
		14'b10110110001001:	sigmoid = 21'b000000000000011001101;
		14'b10110110001010:	sigmoid = 21'b000000000000011001101;
		14'b10110110001011:	sigmoid = 21'b000000000000011001101;
		14'b10110110001100:	sigmoid = 21'b000000000000011001110;
		14'b10110110001101:	sigmoid = 21'b000000000000011001110;
		14'b10110110001110:	sigmoid = 21'b000000000000011001111;
		14'b10110110001111:	sigmoid = 21'b000000000000011001111;
		14'b10110110010000:	sigmoid = 21'b000000000000011001111;
		14'b10110110010001:	sigmoid = 21'b000000000000011010000;
		14'b10110110010010:	sigmoid = 21'b000000000000011010000;
		14'b10110110010011:	sigmoid = 21'b000000000000011010001;
		14'b10110110010100:	sigmoid = 21'b000000000000011010001;
		14'b10110110010101:	sigmoid = 21'b000000000000011010001;
		14'b10110110010110:	sigmoid = 21'b000000000000011010010;
		14'b10110110010111:	sigmoid = 21'b000000000000011010010;
		14'b10110110011000:	sigmoid = 21'b000000000000011010011;
		14'b10110110011001:	sigmoid = 21'b000000000000011010011;
		14'b10110110011010:	sigmoid = 21'b000000000000011010100;
		14'b10110110011011:	sigmoid = 21'b000000000000011010100;
		14'b10110110011100:	sigmoid = 21'b000000000000011010100;
		14'b10110110011101:	sigmoid = 21'b000000000000011010101;
		14'b10110110011110:	sigmoid = 21'b000000000000011010101;
		14'b10110110011111:	sigmoid = 21'b000000000000011010110;
		14'b10110110100000:	sigmoid = 21'b000000000000011010110;
		14'b10110110100001:	sigmoid = 21'b000000000000011010110;
		14'b10110110100010:	sigmoid = 21'b000000000000011010111;
		14'b10110110100011:	sigmoid = 21'b000000000000011010111;
		14'b10110110100100:	sigmoid = 21'b000000000000011011000;
		14'b10110110100101:	sigmoid = 21'b000000000000011011000;
		14'b10110110100110:	sigmoid = 21'b000000000000011011001;
		14'b10110110100111:	sigmoid = 21'b000000000000011011001;
		14'b10110110101000:	sigmoid = 21'b000000000000011011001;
		14'b10110110101001:	sigmoid = 21'b000000000000011011010;
		14'b10110110101010:	sigmoid = 21'b000000000000011011010;
		14'b10110110101011:	sigmoid = 21'b000000000000011011011;
		14'b10110110101100:	sigmoid = 21'b000000000000011011011;
		14'b10110110101101:	sigmoid = 21'b000000000000011011100;
		14'b10110110101110:	sigmoid = 21'b000000000000011011100;
		14'b10110110101111:	sigmoid = 21'b000000000000011011100;
		14'b10110110110000:	sigmoid = 21'b000000000000011011101;
		14'b10110110110001:	sigmoid = 21'b000000000000011011101;
		14'b10110110110010:	sigmoid = 21'b000000000000011011110;
		14'b10110110110011:	sigmoid = 21'b000000000000011011110;
		14'b10110110110100:	sigmoid = 21'b000000000000011011111;
		14'b10110110110101:	sigmoid = 21'b000000000000011011111;
		14'b10110110110110:	sigmoid = 21'b000000000000011011111;
		14'b10110110110111:	sigmoid = 21'b000000000000011100000;
		14'b10110110111000:	sigmoid = 21'b000000000000011100000;
		14'b10110110111001:	sigmoid = 21'b000000000000011100001;
		14'b10110110111010:	sigmoid = 21'b000000000000011100001;
		14'b10110110111011:	sigmoid = 21'b000000000000011100010;
		14'b10110110111100:	sigmoid = 21'b000000000000011100010;
		14'b10110110111101:	sigmoid = 21'b000000000000011100011;
		14'b10110110111110:	sigmoid = 21'b000000000000011100011;
		14'b10110110111111:	sigmoid = 21'b000000000000011100011;
		14'b10110111000000:	sigmoid = 21'b000000000000011100100;
		14'b10110111000001:	sigmoid = 21'b000000000000011100100;
		14'b10110111000010:	sigmoid = 21'b000000000000011100101;
		14'b10110111000011:	sigmoid = 21'b000000000000011100101;
		14'b10110111000100:	sigmoid = 21'b000000000000011100110;
		14'b10110111000101:	sigmoid = 21'b000000000000011100110;
		14'b10110111000110:	sigmoid = 21'b000000000000011100111;
		14'b10110111000111:	sigmoid = 21'b000000000000011100111;
		14'b10110111001000:	sigmoid = 21'b000000000000011100111;
		14'b10110111001001:	sigmoid = 21'b000000000000011101000;
		14'b10110111001010:	sigmoid = 21'b000000000000011101000;
		14'b10110111001011:	sigmoid = 21'b000000000000011101001;
		14'b10110111001100:	sigmoid = 21'b000000000000011101001;
		14'b10110111001101:	sigmoid = 21'b000000000000011101010;
		14'b10110111001110:	sigmoid = 21'b000000000000011101010;
		14'b10110111001111:	sigmoid = 21'b000000000000011101011;
		14'b10110111010000:	sigmoid = 21'b000000000000011101011;
		14'b10110111010001:	sigmoid = 21'b000000000000011101100;
		14'b10110111010010:	sigmoid = 21'b000000000000011101100;
		14'b10110111010011:	sigmoid = 21'b000000000000011101101;
		14'b10110111010100:	sigmoid = 21'b000000000000011101101;
		14'b10110111010101:	sigmoid = 21'b000000000000011101101;
		14'b10110111010110:	sigmoid = 21'b000000000000011101110;
		14'b10110111010111:	sigmoid = 21'b000000000000011101110;
		14'b10110111011000:	sigmoid = 21'b000000000000011101111;
		14'b10110111011001:	sigmoid = 21'b000000000000011101111;
		14'b10110111011010:	sigmoid = 21'b000000000000011110000;
		14'b10110111011011:	sigmoid = 21'b000000000000011110000;
		14'b10110111011100:	sigmoid = 21'b000000000000011110001;
		14'b10110111011101:	sigmoid = 21'b000000000000011110001;
		14'b10110111011110:	sigmoid = 21'b000000000000011110010;
		14'b10110111011111:	sigmoid = 21'b000000000000011110010;
		14'b10110111100000:	sigmoid = 21'b000000000000011110011;
		14'b10110111100001:	sigmoid = 21'b000000000000011110011;
		14'b10110111100010:	sigmoid = 21'b000000000000011110100;
		14'b10110111100011:	sigmoid = 21'b000000000000011110100;
		14'b10110111100100:	sigmoid = 21'b000000000000011110101;
		14'b10110111100101:	sigmoid = 21'b000000000000011110101;
		14'b10110111100110:	sigmoid = 21'b000000000000011110101;
		14'b10110111100111:	sigmoid = 21'b000000000000011110110;
		14'b10110111101000:	sigmoid = 21'b000000000000011110110;
		14'b10110111101001:	sigmoid = 21'b000000000000011110111;
		14'b10110111101010:	sigmoid = 21'b000000000000011110111;
		14'b10110111101011:	sigmoid = 21'b000000000000011111000;
		14'b10110111101100:	sigmoid = 21'b000000000000011111000;
		14'b10110111101101:	sigmoid = 21'b000000000000011111001;
		14'b10110111101110:	sigmoid = 21'b000000000000011111001;
		14'b10110111101111:	sigmoid = 21'b000000000000011111010;
		14'b10110111110000:	sigmoid = 21'b000000000000011111010;
		14'b10110111110001:	sigmoid = 21'b000000000000011111011;
		14'b10110111110010:	sigmoid = 21'b000000000000011111011;
		14'b10110111110011:	sigmoid = 21'b000000000000011111100;
		14'b10110111110100:	sigmoid = 21'b000000000000011111100;
		14'b10110111110101:	sigmoid = 21'b000000000000011111101;
		14'b10110111110110:	sigmoid = 21'b000000000000011111101;
		14'b10110111110111:	sigmoid = 21'b000000000000011111110;
		14'b10110111111000:	sigmoid = 21'b000000000000011111110;
		14'b10110111111001:	sigmoid = 21'b000000000000011111111;
		14'b10110111111010:	sigmoid = 21'b000000000000011111111;
		14'b10110111111011:	sigmoid = 21'b000000000000100000000;
		14'b10110111111100:	sigmoid = 21'b000000000000100000000;
		14'b10110111111101:	sigmoid = 21'b000000000000100000001;
		14'b10110111111110:	sigmoid = 21'b000000000000100000001;
		14'b10110111111111:	sigmoid = 21'b000000000000100000010;
		14'b10111000000000:	sigmoid = 21'b000000000000100000010;
		14'b10111000000001:	sigmoid = 21'b000000000000100000011;
		14'b10111000000010:	sigmoid = 21'b000000000000100000011;
		14'b10111000000011:	sigmoid = 21'b000000000000100000100;
		14'b10111000000100:	sigmoid = 21'b000000000000100000100;
		14'b10111000000101:	sigmoid = 21'b000000000000100000101;
		14'b10111000000110:	sigmoid = 21'b000000000000100000101;
		14'b10111000000111:	sigmoid = 21'b000000000000100000110;
		14'b10111000001000:	sigmoid = 21'b000000000000100000110;
		14'b10111000001001:	sigmoid = 21'b000000000000100000111;
		14'b10111000001010:	sigmoid = 21'b000000000000100000111;
		14'b10111000001011:	sigmoid = 21'b000000000000100001000;
		14'b10111000001100:	sigmoid = 21'b000000000000100001000;
		14'b10111000001101:	sigmoid = 21'b000000000000100001001;
		14'b10111000001110:	sigmoid = 21'b000000000000100001001;
		14'b10111000001111:	sigmoid = 21'b000000000000100001010;
		14'b10111000010000:	sigmoid = 21'b000000000000100001010;
		14'b10111000010001:	sigmoid = 21'b000000000000100001011;
		14'b10111000010010:	sigmoid = 21'b000000000000100001100;
		14'b10111000010011:	sigmoid = 21'b000000000000100001100;
		14'b10111000010100:	sigmoid = 21'b000000000000100001101;
		14'b10111000010101:	sigmoid = 21'b000000000000100001101;
		14'b10111000010110:	sigmoid = 21'b000000000000100001110;
		14'b10111000010111:	sigmoid = 21'b000000000000100001110;
		14'b10111000011000:	sigmoid = 21'b000000000000100001111;
		14'b10111000011001:	sigmoid = 21'b000000000000100001111;
		14'b10111000011010:	sigmoid = 21'b000000000000100010000;
		14'b10111000011011:	sigmoid = 21'b000000000000100010000;
		14'b10111000011100:	sigmoid = 21'b000000000000100010001;
		14'b10111000011101:	sigmoid = 21'b000000000000100010001;
		14'b10111000011110:	sigmoid = 21'b000000000000100010010;
		14'b10111000011111:	sigmoid = 21'b000000000000100010010;
		14'b10111000100000:	sigmoid = 21'b000000000000100010011;
		14'b10111000100001:	sigmoid = 21'b000000000000100010100;
		14'b10111000100010:	sigmoid = 21'b000000000000100010100;
		14'b10111000100011:	sigmoid = 21'b000000000000100010101;
		14'b10111000100100:	sigmoid = 21'b000000000000100010101;
		14'b10111000100101:	sigmoid = 21'b000000000000100010110;
		14'b10111000100110:	sigmoid = 21'b000000000000100010110;
		14'b10111000100111:	sigmoid = 21'b000000000000100010111;
		14'b10111000101000:	sigmoid = 21'b000000000000100010111;
		14'b10111000101001:	sigmoid = 21'b000000000000100011000;
		14'b10111000101010:	sigmoid = 21'b000000000000100011000;
		14'b10111000101011:	sigmoid = 21'b000000000000100011001;
		14'b10111000101100:	sigmoid = 21'b000000000000100011001;
		14'b10111000101101:	sigmoid = 21'b000000000000100011010;
		14'b10111000101110:	sigmoid = 21'b000000000000100011011;
		14'b10111000101111:	sigmoid = 21'b000000000000100011011;
		14'b10111000110000:	sigmoid = 21'b000000000000100011100;
		14'b10111000110001:	sigmoid = 21'b000000000000100011100;
		14'b10111000110010:	sigmoid = 21'b000000000000100011101;
		14'b10111000110011:	sigmoid = 21'b000000000000100011101;
		14'b10111000110100:	sigmoid = 21'b000000000000100011110;
		14'b10111000110101:	sigmoid = 21'b000000000000100011110;
		14'b10111000110110:	sigmoid = 21'b000000000000100011111;
		14'b10111000110111:	sigmoid = 21'b000000000000100100000;
		14'b10111000111000:	sigmoid = 21'b000000000000100100000;
		14'b10111000111001:	sigmoid = 21'b000000000000100100001;
		14'b10111000111010:	sigmoid = 21'b000000000000100100001;
		14'b10111000111011:	sigmoid = 21'b000000000000100100010;
		14'b10111000111100:	sigmoid = 21'b000000000000100100010;
		14'b10111000111101:	sigmoid = 21'b000000000000100100011;
		14'b10111000111110:	sigmoid = 21'b000000000000100100100;
		14'b10111000111111:	sigmoid = 21'b000000000000100100100;
		14'b10111001000000:	sigmoid = 21'b000000000000100100101;
		14'b10111001000001:	sigmoid = 21'b000000000000100100101;
		14'b10111001000010:	sigmoid = 21'b000000000000100100110;
		14'b10111001000011:	sigmoid = 21'b000000000000100100110;
		14'b10111001000100:	sigmoid = 21'b000000000000100100111;
		14'b10111001000101:	sigmoid = 21'b000000000000100101000;
		14'b10111001000110:	sigmoid = 21'b000000000000100101000;
		14'b10111001000111:	sigmoid = 21'b000000000000100101001;
		14'b10111001001000:	sigmoid = 21'b000000000000100101001;
		14'b10111001001001:	sigmoid = 21'b000000000000100101010;
		14'b10111001001010:	sigmoid = 21'b000000000000100101011;
		14'b10111001001011:	sigmoid = 21'b000000000000100101011;
		14'b10111001001100:	sigmoid = 21'b000000000000100101100;
		14'b10111001001101:	sigmoid = 21'b000000000000100101100;
		14'b10111001001110:	sigmoid = 21'b000000000000100101101;
		14'b10111001001111:	sigmoid = 21'b000000000000100101101;
		14'b10111001010000:	sigmoid = 21'b000000000000100101110;
		14'b10111001010001:	sigmoid = 21'b000000000000100101111;
		14'b10111001010010:	sigmoid = 21'b000000000000100101111;
		14'b10111001010011:	sigmoid = 21'b000000000000100110000;
		14'b10111001010100:	sigmoid = 21'b000000000000100110000;
		14'b10111001010101:	sigmoid = 21'b000000000000100110001;
		14'b10111001010110:	sigmoid = 21'b000000000000100110010;
		14'b10111001010111:	sigmoid = 21'b000000000000100110010;
		14'b10111001011000:	sigmoid = 21'b000000000000100110011;
		14'b10111001011001:	sigmoid = 21'b000000000000100110011;
		14'b10111001011010:	sigmoid = 21'b000000000000100110100;
		14'b10111001011011:	sigmoid = 21'b000000000000100110101;
		14'b10111001011100:	sigmoid = 21'b000000000000100110101;
		14'b10111001011101:	sigmoid = 21'b000000000000100110110;
		14'b10111001011110:	sigmoid = 21'b000000000000100110110;
		14'b10111001011111:	sigmoid = 21'b000000000000100110111;
		14'b10111001100000:	sigmoid = 21'b000000000000100111000;
		14'b10111001100001:	sigmoid = 21'b000000000000100111000;
		14'b10111001100010:	sigmoid = 21'b000000000000100111001;
		14'b10111001100011:	sigmoid = 21'b000000000000100111001;
		14'b10111001100100:	sigmoid = 21'b000000000000100111010;
		14'b10111001100101:	sigmoid = 21'b000000000000100111011;
		14'b10111001100110:	sigmoid = 21'b000000000000100111011;
		14'b10111001100111:	sigmoid = 21'b000000000000100111100;
		14'b10111001101000:	sigmoid = 21'b000000000000100111101;
		14'b10111001101001:	sigmoid = 21'b000000000000100111101;
		14'b10111001101010:	sigmoid = 21'b000000000000100111110;
		14'b10111001101011:	sigmoid = 21'b000000000000100111110;
		14'b10111001101100:	sigmoid = 21'b000000000000100111111;
		14'b10111001101101:	sigmoid = 21'b000000000000101000000;
		14'b10111001101110:	sigmoid = 21'b000000000000101000000;
		14'b10111001101111:	sigmoid = 21'b000000000000101000001;
		14'b10111001110000:	sigmoid = 21'b000000000000101000010;
		14'b10111001110001:	sigmoid = 21'b000000000000101000010;
		14'b10111001110010:	sigmoid = 21'b000000000000101000011;
		14'b10111001110011:	sigmoid = 21'b000000000000101000011;
		14'b10111001110100:	sigmoid = 21'b000000000000101000100;
		14'b10111001110101:	sigmoid = 21'b000000000000101000101;
		14'b10111001110110:	sigmoid = 21'b000000000000101000101;
		14'b10111001110111:	sigmoid = 21'b000000000000101000110;
		14'b10111001111000:	sigmoid = 21'b000000000000101000111;
		14'b10111001111001:	sigmoid = 21'b000000000000101000111;
		14'b10111001111010:	sigmoid = 21'b000000000000101001000;
		14'b10111001111011:	sigmoid = 21'b000000000000101001001;
		14'b10111001111100:	sigmoid = 21'b000000000000101001001;
		14'b10111001111101:	sigmoid = 21'b000000000000101001010;
		14'b10111001111110:	sigmoid = 21'b000000000000101001010;
		14'b10111001111111:	sigmoid = 21'b000000000000101001011;
		14'b10111010000000:	sigmoid = 21'b000000000000101001100;
		14'b10111010000001:	sigmoid = 21'b000000000000101001100;
		14'b10111010000010:	sigmoid = 21'b000000000000101001101;
		14'b10111010000011:	sigmoid = 21'b000000000000101001110;
		14'b10111010000100:	sigmoid = 21'b000000000000101001110;
		14'b10111010000101:	sigmoid = 21'b000000000000101001111;
		14'b10111010000110:	sigmoid = 21'b000000000000101010000;
		14'b10111010000111:	sigmoid = 21'b000000000000101010000;
		14'b10111010001000:	sigmoid = 21'b000000000000101010001;
		14'b10111010001001:	sigmoid = 21'b000000000000101010010;
		14'b10111010001010:	sigmoid = 21'b000000000000101010010;
		14'b10111010001011:	sigmoid = 21'b000000000000101010011;
		14'b10111010001100:	sigmoid = 21'b000000000000101010100;
		14'b10111010001101:	sigmoid = 21'b000000000000101010100;
		14'b10111010001110:	sigmoid = 21'b000000000000101010101;
		14'b10111010001111:	sigmoid = 21'b000000000000101010110;
		14'b10111010010000:	sigmoid = 21'b000000000000101010110;
		14'b10111010010001:	sigmoid = 21'b000000000000101010111;
		14'b10111010010010:	sigmoid = 21'b000000000000101011000;
		14'b10111010010011:	sigmoid = 21'b000000000000101011000;
		14'b10111010010100:	sigmoid = 21'b000000000000101011001;
		14'b10111010010101:	sigmoid = 21'b000000000000101011010;
		14'b10111010010110:	sigmoid = 21'b000000000000101011010;
		14'b10111010010111:	sigmoid = 21'b000000000000101011011;
		14'b10111010011000:	sigmoid = 21'b000000000000101011100;
		14'b10111010011001:	sigmoid = 21'b000000000000101011100;
		14'b10111010011010:	sigmoid = 21'b000000000000101011101;
		14'b10111010011011:	sigmoid = 21'b000000000000101011110;
		14'b10111010011100:	sigmoid = 21'b000000000000101011110;
		14'b10111010011101:	sigmoid = 21'b000000000000101011111;
		14'b10111010011110:	sigmoid = 21'b000000000000101100000;
		14'b10111010011111:	sigmoid = 21'b000000000000101100001;
		14'b10111010100000:	sigmoid = 21'b000000000000101100001;
		14'b10111010100001:	sigmoid = 21'b000000000000101100010;
		14'b10111010100010:	sigmoid = 21'b000000000000101100011;
		14'b10111010100011:	sigmoid = 21'b000000000000101100011;
		14'b10111010100100:	sigmoid = 21'b000000000000101100100;
		14'b10111010100101:	sigmoid = 21'b000000000000101100101;
		14'b10111010100110:	sigmoid = 21'b000000000000101100101;
		14'b10111010100111:	sigmoid = 21'b000000000000101100110;
		14'b10111010101000:	sigmoid = 21'b000000000000101100111;
		14'b10111010101001:	sigmoid = 21'b000000000000101100111;
		14'b10111010101010:	sigmoid = 21'b000000000000101101000;
		14'b10111010101011:	sigmoid = 21'b000000000000101101001;
		14'b10111010101100:	sigmoid = 21'b000000000000101101010;
		14'b10111010101101:	sigmoid = 21'b000000000000101101010;
		14'b10111010101110:	sigmoid = 21'b000000000000101101011;
		14'b10111010101111:	sigmoid = 21'b000000000000101101100;
		14'b10111010110000:	sigmoid = 21'b000000000000101101100;
		14'b10111010110001:	sigmoid = 21'b000000000000101101101;
		14'b10111010110010:	sigmoid = 21'b000000000000101101110;
		14'b10111010110011:	sigmoid = 21'b000000000000101101111;
		14'b10111010110100:	sigmoid = 21'b000000000000101101111;
		14'b10111010110101:	sigmoid = 21'b000000000000101110000;
		14'b10111010110110:	sigmoid = 21'b000000000000101110001;
		14'b10111010110111:	sigmoid = 21'b000000000000101110001;
		14'b10111010111000:	sigmoid = 21'b000000000000101110010;
		14'b10111010111001:	sigmoid = 21'b000000000000101110011;
		14'b10111010111010:	sigmoid = 21'b000000000000101110100;
		14'b10111010111011:	sigmoid = 21'b000000000000101110100;
		14'b10111010111100:	sigmoid = 21'b000000000000101110101;
		14'b10111010111101:	sigmoid = 21'b000000000000101110110;
		14'b10111010111110:	sigmoid = 21'b000000000000101110111;
		14'b10111010111111:	sigmoid = 21'b000000000000101110111;
		14'b10111011000000:	sigmoid = 21'b000000000000101111000;
		14'b10111011000001:	sigmoid = 21'b000000000000101111001;
		14'b10111011000010:	sigmoid = 21'b000000000000101111001;
		14'b10111011000011:	sigmoid = 21'b000000000000101111010;
		14'b10111011000100:	sigmoid = 21'b000000000000101111011;
		14'b10111011000101:	sigmoid = 21'b000000000000101111100;
		14'b10111011000110:	sigmoid = 21'b000000000000101111100;
		14'b10111011000111:	sigmoid = 21'b000000000000101111101;
		14'b10111011001000:	sigmoid = 21'b000000000000101111110;
		14'b10111011001001:	sigmoid = 21'b000000000000101111111;
		14'b10111011001010:	sigmoid = 21'b000000000000101111111;
		14'b10111011001011:	sigmoid = 21'b000000000000110000000;
		14'b10111011001100:	sigmoid = 21'b000000000000110000001;
		14'b10111011001101:	sigmoid = 21'b000000000000110000010;
		14'b10111011001110:	sigmoid = 21'b000000000000110000010;
		14'b10111011001111:	sigmoid = 21'b000000000000110000011;
		14'b10111011010000:	sigmoid = 21'b000000000000110000100;
		14'b10111011010001:	sigmoid = 21'b000000000000110000101;
		14'b10111011010010:	sigmoid = 21'b000000000000110000101;
		14'b10111011010011:	sigmoid = 21'b000000000000110000110;
		14'b10111011010100:	sigmoid = 21'b000000000000110000111;
		14'b10111011010101:	sigmoid = 21'b000000000000110001000;
		14'b10111011010110:	sigmoid = 21'b000000000000110001001;
		14'b10111011010111:	sigmoid = 21'b000000000000110001001;
		14'b10111011011000:	sigmoid = 21'b000000000000110001010;
		14'b10111011011001:	sigmoid = 21'b000000000000110001011;
		14'b10111011011010:	sigmoid = 21'b000000000000110001100;
		14'b10111011011011:	sigmoid = 21'b000000000000110001100;
		14'b10111011011100:	sigmoid = 21'b000000000000110001101;
		14'b10111011011101:	sigmoid = 21'b000000000000110001110;
		14'b10111011011110:	sigmoid = 21'b000000000000110001111;
		14'b10111011011111:	sigmoid = 21'b000000000000110001111;
		14'b10111011100000:	sigmoid = 21'b000000000000110010000;
		14'b10111011100001:	sigmoid = 21'b000000000000110010001;
		14'b10111011100010:	sigmoid = 21'b000000000000110010010;
		14'b10111011100011:	sigmoid = 21'b000000000000110010011;
		14'b10111011100100:	sigmoid = 21'b000000000000110010011;
		14'b10111011100101:	sigmoid = 21'b000000000000110010100;
		14'b10111011100110:	sigmoid = 21'b000000000000110010101;
		14'b10111011100111:	sigmoid = 21'b000000000000110010110;
		14'b10111011101000:	sigmoid = 21'b000000000000110010111;
		14'b10111011101001:	sigmoid = 21'b000000000000110010111;
		14'b10111011101010:	sigmoid = 21'b000000000000110011000;
		14'b10111011101011:	sigmoid = 21'b000000000000110011001;
		14'b10111011101100:	sigmoid = 21'b000000000000110011010;
		14'b10111011101101:	sigmoid = 21'b000000000000110011011;
		14'b10111011101110:	sigmoid = 21'b000000000000110011011;
		14'b10111011101111:	sigmoid = 21'b000000000000110011100;
		14'b10111011110000:	sigmoid = 21'b000000000000110011101;
		14'b10111011110001:	sigmoid = 21'b000000000000110011110;
		14'b10111011110010:	sigmoid = 21'b000000000000110011111;
		14'b10111011110011:	sigmoid = 21'b000000000000110011111;
		14'b10111011110100:	sigmoid = 21'b000000000000110100000;
		14'b10111011110101:	sigmoid = 21'b000000000000110100001;
		14'b10111011110110:	sigmoid = 21'b000000000000110100010;
		14'b10111011110111:	sigmoid = 21'b000000000000110100011;
		14'b10111011111000:	sigmoid = 21'b000000000000110100100;
		14'b10111011111001:	sigmoid = 21'b000000000000110100100;
		14'b10111011111010:	sigmoid = 21'b000000000000110100101;
		14'b10111011111011:	sigmoid = 21'b000000000000110100110;
		14'b10111011111100:	sigmoid = 21'b000000000000110100111;
		14'b10111011111101:	sigmoid = 21'b000000000000110101000;
		14'b10111011111110:	sigmoid = 21'b000000000000110101000;
		14'b10111011111111:	sigmoid = 21'b000000000000110101001;
		14'b10111100000000:	sigmoid = 21'b000000000000110101010;
		14'b10111100000001:	sigmoid = 21'b000000000000110101011;
		14'b10111100000010:	sigmoid = 21'b000000000000110101100;
		14'b10111100000011:	sigmoid = 21'b000000000000110101101;
		14'b10111100000100:	sigmoid = 21'b000000000000110101101;
		14'b10111100000101:	sigmoid = 21'b000000000000110101110;
		14'b10111100000110:	sigmoid = 21'b000000000000110101111;
		14'b10111100000111:	sigmoid = 21'b000000000000110110000;
		14'b10111100001000:	sigmoid = 21'b000000000000110110001;
		14'b10111100001001:	sigmoid = 21'b000000000000110110010;
		14'b10111100001010:	sigmoid = 21'b000000000000110110011;
		14'b10111100001011:	sigmoid = 21'b000000000000110110011;
		14'b10111100001100:	sigmoid = 21'b000000000000110110100;
		14'b10111100001101:	sigmoid = 21'b000000000000110110101;
		14'b10111100001110:	sigmoid = 21'b000000000000110110110;
		14'b10111100001111:	sigmoid = 21'b000000000000110110111;
		14'b10111100010000:	sigmoid = 21'b000000000000110111000;
		14'b10111100010001:	sigmoid = 21'b000000000000110111001;
		14'b10111100010010:	sigmoid = 21'b000000000000110111001;
		14'b10111100010011:	sigmoid = 21'b000000000000110111010;
		14'b10111100010100:	sigmoid = 21'b000000000000110111011;
		14'b10111100010101:	sigmoid = 21'b000000000000110111100;
		14'b10111100010110:	sigmoid = 21'b000000000000110111101;
		14'b10111100010111:	sigmoid = 21'b000000000000110111110;
		14'b10111100011000:	sigmoid = 21'b000000000000110111111;
		14'b10111100011001:	sigmoid = 21'b000000000000110111111;
		14'b10111100011010:	sigmoid = 21'b000000000000111000000;
		14'b10111100011011:	sigmoid = 21'b000000000000111000001;
		14'b10111100011100:	sigmoid = 21'b000000000000111000010;
		14'b10111100011101:	sigmoid = 21'b000000000000111000011;
		14'b10111100011110:	sigmoid = 21'b000000000000111000100;
		14'b10111100011111:	sigmoid = 21'b000000000000111000101;
		14'b10111100100000:	sigmoid = 21'b000000000000111000110;
		14'b10111100100001:	sigmoid = 21'b000000000000111000111;
		14'b10111100100010:	sigmoid = 21'b000000000000111000111;
		14'b10111100100011:	sigmoid = 21'b000000000000111001000;
		14'b10111100100100:	sigmoid = 21'b000000000000111001001;
		14'b10111100100101:	sigmoid = 21'b000000000000111001010;
		14'b10111100100110:	sigmoid = 21'b000000000000111001011;
		14'b10111100100111:	sigmoid = 21'b000000000000111001100;
		14'b10111100101000:	sigmoid = 21'b000000000000111001101;
		14'b10111100101001:	sigmoid = 21'b000000000000111001110;
		14'b10111100101010:	sigmoid = 21'b000000000000111001111;
		14'b10111100101011:	sigmoid = 21'b000000000000111001111;
		14'b10111100101100:	sigmoid = 21'b000000000000111010000;
		14'b10111100101101:	sigmoid = 21'b000000000000111010001;
		14'b10111100101110:	sigmoid = 21'b000000000000111010010;
		14'b10111100101111:	sigmoid = 21'b000000000000111010011;
		14'b10111100110000:	sigmoid = 21'b000000000000111010100;
		14'b10111100110001:	sigmoid = 21'b000000000000111010101;
		14'b10111100110010:	sigmoid = 21'b000000000000111010110;
		14'b10111100110011:	sigmoid = 21'b000000000000111010111;
		14'b10111100110100:	sigmoid = 21'b000000000000111011000;
		14'b10111100110101:	sigmoid = 21'b000000000000111011001;
		14'b10111100110110:	sigmoid = 21'b000000000000111011010;
		14'b10111100110111:	sigmoid = 21'b000000000000111011010;
		14'b10111100111000:	sigmoid = 21'b000000000000111011011;
		14'b10111100111001:	sigmoid = 21'b000000000000111011100;
		14'b10111100111010:	sigmoid = 21'b000000000000111011101;
		14'b10111100111011:	sigmoid = 21'b000000000000111011110;
		14'b10111100111100:	sigmoid = 21'b000000000000111011111;
		14'b10111100111101:	sigmoid = 21'b000000000000111100000;
		14'b10111100111110:	sigmoid = 21'b000000000000111100001;
		14'b10111100111111:	sigmoid = 21'b000000000000111100010;
		14'b10111101000000:	sigmoid = 21'b000000000000111100011;
		14'b10111101000001:	sigmoid = 21'b000000000000111100100;
		14'b10111101000010:	sigmoid = 21'b000000000000111100101;
		14'b10111101000011:	sigmoid = 21'b000000000000111100110;
		14'b10111101000100:	sigmoid = 21'b000000000000111100111;
		14'b10111101000101:	sigmoid = 21'b000000000000111101000;
		14'b10111101000110:	sigmoid = 21'b000000000000111101001;
		14'b10111101000111:	sigmoid = 21'b000000000000111101010;
		14'b10111101001000:	sigmoid = 21'b000000000000111101011;
		14'b10111101001001:	sigmoid = 21'b000000000000111101011;
		14'b10111101001010:	sigmoid = 21'b000000000000111101100;
		14'b10111101001011:	sigmoid = 21'b000000000000111101101;
		14'b10111101001100:	sigmoid = 21'b000000000000111101110;
		14'b10111101001101:	sigmoid = 21'b000000000000111101111;
		14'b10111101001110:	sigmoid = 21'b000000000000111110000;
		14'b10111101001111:	sigmoid = 21'b000000000000111110001;
		14'b10111101010000:	sigmoid = 21'b000000000000111110010;
		14'b10111101010001:	sigmoid = 21'b000000000000111110011;
		14'b10111101010010:	sigmoid = 21'b000000000000111110100;
		14'b10111101010011:	sigmoid = 21'b000000000000111110101;
		14'b10111101010100:	sigmoid = 21'b000000000000111110110;
		14'b10111101010101:	sigmoid = 21'b000000000000111110111;
		14'b10111101010110:	sigmoid = 21'b000000000000111111000;
		14'b10111101010111:	sigmoid = 21'b000000000000111111001;
		14'b10111101011000:	sigmoid = 21'b000000000000111111010;
		14'b10111101011001:	sigmoid = 21'b000000000000111111011;
		14'b10111101011010:	sigmoid = 21'b000000000000111111100;
		14'b10111101011011:	sigmoid = 21'b000000000000111111101;
		14'b10111101011100:	sigmoid = 21'b000000000000111111110;
		14'b10111101011101:	sigmoid = 21'b000000000000111111111;
		14'b10111101011110:	sigmoid = 21'b000000000001000000000;
		14'b10111101011111:	sigmoid = 21'b000000000001000000001;
		14'b10111101100000:	sigmoid = 21'b000000000001000000010;
		14'b10111101100001:	sigmoid = 21'b000000000001000000011;
		14'b10111101100010:	sigmoid = 21'b000000000001000000100;
		14'b10111101100011:	sigmoid = 21'b000000000001000000101;
		14'b10111101100100:	sigmoid = 21'b000000000001000000110;
		14'b10111101100101:	sigmoid = 21'b000000000001000000111;
		14'b10111101100110:	sigmoid = 21'b000000000001000001000;
		14'b10111101100111:	sigmoid = 21'b000000000001000001001;
		14'b10111101101000:	sigmoid = 21'b000000000001000001010;
		14'b10111101101001:	sigmoid = 21'b000000000001000001011;
		14'b10111101101010:	sigmoid = 21'b000000000001000001100;
		14'b10111101101011:	sigmoid = 21'b000000000001000001101;
		14'b10111101101100:	sigmoid = 21'b000000000001000001110;
		14'b10111101101101:	sigmoid = 21'b000000000001000001111;
		14'b10111101101110:	sigmoid = 21'b000000000001000010000;
		14'b10111101101111:	sigmoid = 21'b000000000001000010001;
		14'b10111101110000:	sigmoid = 21'b000000000001000010010;
		14'b10111101110001:	sigmoid = 21'b000000000001000010011;
		14'b10111101110010:	sigmoid = 21'b000000000001000010100;
		14'b10111101110011:	sigmoid = 21'b000000000001000010110;
		14'b10111101110100:	sigmoid = 21'b000000000001000010111;
		14'b10111101110101:	sigmoid = 21'b000000000001000011000;
		14'b10111101110110:	sigmoid = 21'b000000000001000011001;
		14'b10111101110111:	sigmoid = 21'b000000000001000011010;
		14'b10111101111000:	sigmoid = 21'b000000000001000011011;
		14'b10111101111001:	sigmoid = 21'b000000000001000011100;
		14'b10111101111010:	sigmoid = 21'b000000000001000011101;
		14'b10111101111011:	sigmoid = 21'b000000000001000011110;
		14'b10111101111100:	sigmoid = 21'b000000000001000011111;
		14'b10111101111101:	sigmoid = 21'b000000000001000100000;
		14'b10111101111110:	sigmoid = 21'b000000000001000100001;
		14'b10111101111111:	sigmoid = 21'b000000000001000100010;
		14'b10111110000000:	sigmoid = 21'b000000000001000100011;
		14'b10111110000001:	sigmoid = 21'b000000000001000100100;
		14'b10111110000010:	sigmoid = 21'b000000000001000100101;
		14'b10111110000011:	sigmoid = 21'b000000000001000100110;
		14'b10111110000100:	sigmoid = 21'b000000000001000101000;
		14'b10111110000101:	sigmoid = 21'b000000000001000101001;
		14'b10111110000110:	sigmoid = 21'b000000000001000101010;
		14'b10111110000111:	sigmoid = 21'b000000000001000101011;
		14'b10111110001000:	sigmoid = 21'b000000000001000101100;
		14'b10111110001001:	sigmoid = 21'b000000000001000101101;
		14'b10111110001010:	sigmoid = 21'b000000000001000101110;
		14'b10111110001011:	sigmoid = 21'b000000000001000101111;
		14'b10111110001100:	sigmoid = 21'b000000000001000110000;
		14'b10111110001101:	sigmoid = 21'b000000000001000110001;
		14'b10111110001110:	sigmoid = 21'b000000000001000110010;
		14'b10111110001111:	sigmoid = 21'b000000000001000110100;
		14'b10111110010000:	sigmoid = 21'b000000000001000110101;
		14'b10111110010001:	sigmoid = 21'b000000000001000110110;
		14'b10111110010010:	sigmoid = 21'b000000000001000110111;
		14'b10111110010011:	sigmoid = 21'b000000000001000111000;
		14'b10111110010100:	sigmoid = 21'b000000000001000111001;
		14'b10111110010101:	sigmoid = 21'b000000000001000111010;
		14'b10111110010110:	sigmoid = 21'b000000000001000111011;
		14'b10111110010111:	sigmoid = 21'b000000000001000111100;
		14'b10111110011000:	sigmoid = 21'b000000000001000111110;
		14'b10111110011001:	sigmoid = 21'b000000000001000111111;
		14'b10111110011010:	sigmoid = 21'b000000000001001000000;
		14'b10111110011011:	sigmoid = 21'b000000000001001000001;
		14'b10111110011100:	sigmoid = 21'b000000000001001000010;
		14'b10111110011101:	sigmoid = 21'b000000000001001000011;
		14'b10111110011110:	sigmoid = 21'b000000000001001000100;
		14'b10111110011111:	sigmoid = 21'b000000000001001000101;
		14'b10111110100000:	sigmoid = 21'b000000000001001000111;
		14'b10111110100001:	sigmoid = 21'b000000000001001001000;
		14'b10111110100010:	sigmoid = 21'b000000000001001001001;
		14'b10111110100011:	sigmoid = 21'b000000000001001001010;
		14'b10111110100100:	sigmoid = 21'b000000000001001001011;
		14'b10111110100101:	sigmoid = 21'b000000000001001001100;
		14'b10111110100110:	sigmoid = 21'b000000000001001001101;
		14'b10111110100111:	sigmoid = 21'b000000000001001001111;
		14'b10111110101000:	sigmoid = 21'b000000000001001010000;
		14'b10111110101001:	sigmoid = 21'b000000000001001010001;
		14'b10111110101010:	sigmoid = 21'b000000000001001010010;
		14'b10111110101011:	sigmoid = 21'b000000000001001010011;
		14'b10111110101100:	sigmoid = 21'b000000000001001010100;
		14'b10111110101101:	sigmoid = 21'b000000000001001010110;
		14'b10111110101110:	sigmoid = 21'b000000000001001010111;
		14'b10111110101111:	sigmoid = 21'b000000000001001011000;
		14'b10111110110000:	sigmoid = 21'b000000000001001011001;
		14'b10111110110001:	sigmoid = 21'b000000000001001011010;
		14'b10111110110010:	sigmoid = 21'b000000000001001011011;
		14'b10111110110011:	sigmoid = 21'b000000000001001011101;
		14'b10111110110100:	sigmoid = 21'b000000000001001011110;
		14'b10111110110101:	sigmoid = 21'b000000000001001011111;
		14'b10111110110110:	sigmoid = 21'b000000000001001100000;
		14'b10111110110111:	sigmoid = 21'b000000000001001100001;
		14'b10111110111000:	sigmoid = 21'b000000000001001100011;
		14'b10111110111001:	sigmoid = 21'b000000000001001100100;
		14'b10111110111010:	sigmoid = 21'b000000000001001100101;
		14'b10111110111011:	sigmoid = 21'b000000000001001100110;
		14'b10111110111100:	sigmoid = 21'b000000000001001100111;
		14'b10111110111101:	sigmoid = 21'b000000000001001101001;
		14'b10111110111110:	sigmoid = 21'b000000000001001101010;
		14'b10111110111111:	sigmoid = 21'b000000000001001101011;
		14'b10111111000000:	sigmoid = 21'b000000000001001101100;
		14'b10111111000001:	sigmoid = 21'b000000000001001101101;
		14'b10111111000010:	sigmoid = 21'b000000000001001101111;
		14'b10111111000011:	sigmoid = 21'b000000000001001110000;
		14'b10111111000100:	sigmoid = 21'b000000000001001110001;
		14'b10111111000101:	sigmoid = 21'b000000000001001110010;
		14'b10111111000110:	sigmoid = 21'b000000000001001110011;
		14'b10111111000111:	sigmoid = 21'b000000000001001110101;
		14'b10111111001000:	sigmoid = 21'b000000000001001110110;
		14'b10111111001001:	sigmoid = 21'b000000000001001110111;
		14'b10111111001010:	sigmoid = 21'b000000000001001111000;
		14'b10111111001011:	sigmoid = 21'b000000000001001111010;
		14'b10111111001100:	sigmoid = 21'b000000000001001111011;
		14'b10111111001101:	sigmoid = 21'b000000000001001111100;
		14'b10111111001110:	sigmoid = 21'b000000000001001111101;
		14'b10111111001111:	sigmoid = 21'b000000000001001111111;
		14'b10111111010000:	sigmoid = 21'b000000000001010000000;
		14'b10111111010001:	sigmoid = 21'b000000000001010000001;
		14'b10111111010010:	sigmoid = 21'b000000000001010000010;
		14'b10111111010011:	sigmoid = 21'b000000000001010000100;
		14'b10111111010100:	sigmoid = 21'b000000000001010000101;
		14'b10111111010101:	sigmoid = 21'b000000000001010000110;
		14'b10111111010110:	sigmoid = 21'b000000000001010000111;
		14'b10111111010111:	sigmoid = 21'b000000000001010001001;
		14'b10111111011000:	sigmoid = 21'b000000000001010001010;
		14'b10111111011001:	sigmoid = 21'b000000000001010001011;
		14'b10111111011010:	sigmoid = 21'b000000000001010001100;
		14'b10111111011011:	sigmoid = 21'b000000000001010001110;
		14'b10111111011100:	sigmoid = 21'b000000000001010001111;
		14'b10111111011101:	sigmoid = 21'b000000000001010010000;
		14'b10111111011110:	sigmoid = 21'b000000000001010010010;
		14'b10111111011111:	sigmoid = 21'b000000000001010010011;
		14'b10111111100000:	sigmoid = 21'b000000000001010010100;
		14'b10111111100001:	sigmoid = 21'b000000000001010010101;
		14'b10111111100010:	sigmoid = 21'b000000000001010010111;
		14'b10111111100011:	sigmoid = 21'b000000000001010011000;
		14'b10111111100100:	sigmoid = 21'b000000000001010011001;
		14'b10111111100101:	sigmoid = 21'b000000000001010011011;
		14'b10111111100110:	sigmoid = 21'b000000000001010011100;
		14'b10111111100111:	sigmoid = 21'b000000000001010011101;
		14'b10111111101000:	sigmoid = 21'b000000000001010011111;
		14'b10111111101001:	sigmoid = 21'b000000000001010100000;
		14'b10111111101010:	sigmoid = 21'b000000000001010100001;
		14'b10111111101011:	sigmoid = 21'b000000000001010100011;
		14'b10111111101100:	sigmoid = 21'b000000000001010100100;
		14'b10111111101101:	sigmoid = 21'b000000000001010100101;
		14'b10111111101110:	sigmoid = 21'b000000000001010100110;
		14'b10111111101111:	sigmoid = 21'b000000000001010101000;
		14'b10111111110000:	sigmoid = 21'b000000000001010101001;
		14'b10111111110001:	sigmoid = 21'b000000000001010101010;
		14'b10111111110010:	sigmoid = 21'b000000000001010101100;
		14'b10111111110011:	sigmoid = 21'b000000000001010101101;
		14'b10111111110100:	sigmoid = 21'b000000000001010101110;
		14'b10111111110101:	sigmoid = 21'b000000000001010110000;
		14'b10111111110110:	sigmoid = 21'b000000000001010110001;
		14'b10111111110111:	sigmoid = 21'b000000000001010110011;
		14'b10111111111000:	sigmoid = 21'b000000000001010110100;
		14'b10111111111001:	sigmoid = 21'b000000000001010110101;
		14'b10111111111010:	sigmoid = 21'b000000000001010110111;
		14'b10111111111011:	sigmoid = 21'b000000000001010111000;
		14'b10111111111100:	sigmoid = 21'b000000000001010111001;
		14'b10111111111101:	sigmoid = 21'b000000000001010111011;
		14'b10111111111110:	sigmoid = 21'b000000000001010111100;
		14'b10111111111111:	sigmoid = 21'b000000000001010111101;
		14'b11000000000000:	sigmoid = 21'b000000000001010111111;
		14'b11000000000001:	sigmoid = 21'b000000000001011000000;
		14'b11000000000010:	sigmoid = 21'b000000000001011000010;
		14'b11000000000011:	sigmoid = 21'b000000000001011000011;
		14'b11000000000100:	sigmoid = 21'b000000000001011000100;
		14'b11000000000101:	sigmoid = 21'b000000000001011000110;
		14'b11000000000110:	sigmoid = 21'b000000000001011000111;
		14'b11000000000111:	sigmoid = 21'b000000000001011001000;
		14'b11000000001000:	sigmoid = 21'b000000000001011001010;
		14'b11000000001001:	sigmoid = 21'b000000000001011001011;
		14'b11000000001010:	sigmoid = 21'b000000000001011001101;
		14'b11000000001011:	sigmoid = 21'b000000000001011001110;
		14'b11000000001100:	sigmoid = 21'b000000000001011001111;
		14'b11000000001101:	sigmoid = 21'b000000000001011010001;
		14'b11000000001110:	sigmoid = 21'b000000000001011010010;
		14'b11000000001111:	sigmoid = 21'b000000000001011010100;
		14'b11000000010000:	sigmoid = 21'b000000000001011010101;
		14'b11000000010001:	sigmoid = 21'b000000000001011010111;
		14'b11000000010010:	sigmoid = 21'b000000000001011011000;
		14'b11000000010011:	sigmoid = 21'b000000000001011011001;
		14'b11000000010100:	sigmoid = 21'b000000000001011011011;
		14'b11000000010101:	sigmoid = 21'b000000000001011011100;
		14'b11000000010110:	sigmoid = 21'b000000000001011011110;
		14'b11000000010111:	sigmoid = 21'b000000000001011011111;
		14'b11000000011000:	sigmoid = 21'b000000000001011100001;
		14'b11000000011001:	sigmoid = 21'b000000000001011100010;
		14'b11000000011010:	sigmoid = 21'b000000000001011100011;
		14'b11000000011011:	sigmoid = 21'b000000000001011100101;
		14'b11000000011100:	sigmoid = 21'b000000000001011100110;
		14'b11000000011101:	sigmoid = 21'b000000000001011101000;
		14'b11000000011110:	sigmoid = 21'b000000000001011101001;
		14'b11000000011111:	sigmoid = 21'b000000000001011101011;
		14'b11000000100000:	sigmoid = 21'b000000000001011101100;
		14'b11000000100001:	sigmoid = 21'b000000000001011101110;
		14'b11000000100010:	sigmoid = 21'b000000000001011101111;
		14'b11000000100011:	sigmoid = 21'b000000000001011110001;
		14'b11000000100100:	sigmoid = 21'b000000000001011110010;
		14'b11000000100101:	sigmoid = 21'b000000000001011110011;
		14'b11000000100110:	sigmoid = 21'b000000000001011110101;
		14'b11000000100111:	sigmoid = 21'b000000000001011110110;
		14'b11000000101000:	sigmoid = 21'b000000000001011111000;
		14'b11000000101001:	sigmoid = 21'b000000000001011111001;
		14'b11000000101010:	sigmoid = 21'b000000000001011111011;
		14'b11000000101011:	sigmoid = 21'b000000000001011111100;
		14'b11000000101100:	sigmoid = 21'b000000000001011111110;
		14'b11000000101101:	sigmoid = 21'b000000000001011111111;
		14'b11000000101110:	sigmoid = 21'b000000000001100000001;
		14'b11000000101111:	sigmoid = 21'b000000000001100000010;
		14'b11000000110000:	sigmoid = 21'b000000000001100000100;
		14'b11000000110001:	sigmoid = 21'b000000000001100000101;
		14'b11000000110010:	sigmoid = 21'b000000000001100000111;
		14'b11000000110011:	sigmoid = 21'b000000000001100001000;
		14'b11000000110100:	sigmoid = 21'b000000000001100001010;
		14'b11000000110101:	sigmoid = 21'b000000000001100001011;
		14'b11000000110110:	sigmoid = 21'b000000000001100001101;
		14'b11000000110111:	sigmoid = 21'b000000000001100001111;
		14'b11000000111000:	sigmoid = 21'b000000000001100010000;
		14'b11000000111001:	sigmoid = 21'b000000000001100010010;
		14'b11000000111010:	sigmoid = 21'b000000000001100010011;
		14'b11000000111011:	sigmoid = 21'b000000000001100010101;
		14'b11000000111100:	sigmoid = 21'b000000000001100010110;
		14'b11000000111101:	sigmoid = 21'b000000000001100011000;
		14'b11000000111110:	sigmoid = 21'b000000000001100011001;
		14'b11000000111111:	sigmoid = 21'b000000000001100011011;
		14'b11000001000000:	sigmoid = 21'b000000000001100011100;
		14'b11000001000001:	sigmoid = 21'b000000000001100011110;
		14'b11000001000010:	sigmoid = 21'b000000000001100100000;
		14'b11000001000011:	sigmoid = 21'b000000000001100100001;
		14'b11000001000100:	sigmoid = 21'b000000000001100100011;
		14'b11000001000101:	sigmoid = 21'b000000000001100100100;
		14'b11000001000110:	sigmoid = 21'b000000000001100100110;
		14'b11000001000111:	sigmoid = 21'b000000000001100100111;
		14'b11000001001000:	sigmoid = 21'b000000000001100101001;
		14'b11000001001001:	sigmoid = 21'b000000000001100101011;
		14'b11000001001010:	sigmoid = 21'b000000000001100101100;
		14'b11000001001011:	sigmoid = 21'b000000000001100101110;
		14'b11000001001100:	sigmoid = 21'b000000000001100101111;
		14'b11000001001101:	sigmoid = 21'b000000000001100110001;
		14'b11000001001110:	sigmoid = 21'b000000000001100110010;
		14'b11000001001111:	sigmoid = 21'b000000000001100110100;
		14'b11000001010000:	sigmoid = 21'b000000000001100110110;
		14'b11000001010001:	sigmoid = 21'b000000000001100110111;
		14'b11000001010010:	sigmoid = 21'b000000000001100111001;
		14'b11000001010011:	sigmoid = 21'b000000000001100111011;
		14'b11000001010100:	sigmoid = 21'b000000000001100111100;
		14'b11000001010101:	sigmoid = 21'b000000000001100111110;
		14'b11000001010110:	sigmoid = 21'b000000000001100111111;
		14'b11000001010111:	sigmoid = 21'b000000000001101000001;
		14'b11000001011000:	sigmoid = 21'b000000000001101000011;
		14'b11000001011001:	sigmoid = 21'b000000000001101000100;
		14'b11000001011010:	sigmoid = 21'b000000000001101000110;
		14'b11000001011011:	sigmoid = 21'b000000000001101001000;
		14'b11000001011100:	sigmoid = 21'b000000000001101001001;
		14'b11000001011101:	sigmoid = 21'b000000000001101001011;
		14'b11000001011110:	sigmoid = 21'b000000000001101001100;
		14'b11000001011111:	sigmoid = 21'b000000000001101001110;
		14'b11000001100000:	sigmoid = 21'b000000000001101010000;
		14'b11000001100001:	sigmoid = 21'b000000000001101010001;
		14'b11000001100010:	sigmoid = 21'b000000000001101010011;
		14'b11000001100011:	sigmoid = 21'b000000000001101010101;
		14'b11000001100100:	sigmoid = 21'b000000000001101010110;
		14'b11000001100101:	sigmoid = 21'b000000000001101011000;
		14'b11000001100110:	sigmoid = 21'b000000000001101011010;
		14'b11000001100111:	sigmoid = 21'b000000000001101011011;
		14'b11000001101000:	sigmoid = 21'b000000000001101011101;
		14'b11000001101001:	sigmoid = 21'b000000000001101011111;
		14'b11000001101010:	sigmoid = 21'b000000000001101100000;
		14'b11000001101011:	sigmoid = 21'b000000000001101100010;
		14'b11000001101100:	sigmoid = 21'b000000000001101100100;
		14'b11000001101101:	sigmoid = 21'b000000000001101100110;
		14'b11000001101110:	sigmoid = 21'b000000000001101100111;
		14'b11000001101111:	sigmoid = 21'b000000000001101101001;
		14'b11000001110000:	sigmoid = 21'b000000000001101101011;
		14'b11000001110001:	sigmoid = 21'b000000000001101101100;
		14'b11000001110010:	sigmoid = 21'b000000000001101101110;
		14'b11000001110011:	sigmoid = 21'b000000000001101110000;
		14'b11000001110100:	sigmoid = 21'b000000000001101110010;
		14'b11000001110101:	sigmoid = 21'b000000000001101110011;
		14'b11000001110110:	sigmoid = 21'b000000000001101110101;
		14'b11000001110111:	sigmoid = 21'b000000000001101110111;
		14'b11000001111000:	sigmoid = 21'b000000000001101111000;
		14'b11000001111001:	sigmoid = 21'b000000000001101111010;
		14'b11000001111010:	sigmoid = 21'b000000000001101111100;
		14'b11000001111011:	sigmoid = 21'b000000000001101111110;
		14'b11000001111100:	sigmoid = 21'b000000000001101111111;
		14'b11000001111101:	sigmoid = 21'b000000000001110000001;
		14'b11000001111110:	sigmoid = 21'b000000000001110000011;
		14'b11000001111111:	sigmoid = 21'b000000000001110000101;
		14'b11000010000000:	sigmoid = 21'b000000000001110000110;
		14'b11000010000001:	sigmoid = 21'b000000000001110001000;
		14'b11000010000010:	sigmoid = 21'b000000000001110001010;
		14'b11000010000011:	sigmoid = 21'b000000000001110001100;
		14'b11000010000100:	sigmoid = 21'b000000000001110001110;
		14'b11000010000101:	sigmoid = 21'b000000000001110001111;
		14'b11000010000110:	sigmoid = 21'b000000000001110010001;
		14'b11000010000111:	sigmoid = 21'b000000000001110010011;
		14'b11000010001000:	sigmoid = 21'b000000000001110010101;
		14'b11000010001001:	sigmoid = 21'b000000000001110010110;
		14'b11000010001010:	sigmoid = 21'b000000000001110011000;
		14'b11000010001011:	sigmoid = 21'b000000000001110011010;
		14'b11000010001100:	sigmoid = 21'b000000000001110011100;
		14'b11000010001101:	sigmoid = 21'b000000000001110011110;
		14'b11000010001110:	sigmoid = 21'b000000000001110011111;
		14'b11000010001111:	sigmoid = 21'b000000000001110100001;
		14'b11000010010000:	sigmoid = 21'b000000000001110100011;
		14'b11000010010001:	sigmoid = 21'b000000000001110100101;
		14'b11000010010010:	sigmoid = 21'b000000000001110100111;
		14'b11000010010011:	sigmoid = 21'b000000000001110101001;
		14'b11000010010100:	sigmoid = 21'b000000000001110101010;
		14'b11000010010101:	sigmoid = 21'b000000000001110101100;
		14'b11000010010110:	sigmoid = 21'b000000000001110101110;
		14'b11000010010111:	sigmoid = 21'b000000000001110110000;
		14'b11000010011000:	sigmoid = 21'b000000000001110110010;
		14'b11000010011001:	sigmoid = 21'b000000000001110110100;
		14'b11000010011010:	sigmoid = 21'b000000000001110110101;
		14'b11000010011011:	sigmoid = 21'b000000000001110110111;
		14'b11000010011100:	sigmoid = 21'b000000000001110111001;
		14'b11000010011101:	sigmoid = 21'b000000000001110111011;
		14'b11000010011110:	sigmoid = 21'b000000000001110111101;
		14'b11000010011111:	sigmoid = 21'b000000000001110111111;
		14'b11000010100000:	sigmoid = 21'b000000000001111000001;
		14'b11000010100001:	sigmoid = 21'b000000000001111000011;
		14'b11000010100010:	sigmoid = 21'b000000000001111000100;
		14'b11000010100011:	sigmoid = 21'b000000000001111000110;
		14'b11000010100100:	sigmoid = 21'b000000000001111001000;
		14'b11000010100101:	sigmoid = 21'b000000000001111001010;
		14'b11000010100110:	sigmoid = 21'b000000000001111001100;
		14'b11000010100111:	sigmoid = 21'b000000000001111001110;
		14'b11000010101000:	sigmoid = 21'b000000000001111010000;
		14'b11000010101001:	sigmoid = 21'b000000000001111010010;
		14'b11000010101010:	sigmoid = 21'b000000000001111010100;
		14'b11000010101011:	sigmoid = 21'b000000000001111010110;
		14'b11000010101100:	sigmoid = 21'b000000000001111010111;
		14'b11000010101101:	sigmoid = 21'b000000000001111011001;
		14'b11000010101110:	sigmoid = 21'b000000000001111011011;
		14'b11000010101111:	sigmoid = 21'b000000000001111011101;
		14'b11000010110000:	sigmoid = 21'b000000000001111011111;
		14'b11000010110001:	sigmoid = 21'b000000000001111100001;
		14'b11000010110010:	sigmoid = 21'b000000000001111100011;
		14'b11000010110011:	sigmoid = 21'b000000000001111100101;
		14'b11000010110100:	sigmoid = 21'b000000000001111100111;
		14'b11000010110101:	sigmoid = 21'b000000000001111101001;
		14'b11000010110110:	sigmoid = 21'b000000000001111101011;
		14'b11000010110111:	sigmoid = 21'b000000000001111101101;
		14'b11000010111000:	sigmoid = 21'b000000000001111101111;
		14'b11000010111001:	sigmoid = 21'b000000000001111110001;
		14'b11000010111010:	sigmoid = 21'b000000000001111110011;
		14'b11000010111011:	sigmoid = 21'b000000000001111110101;
		14'b11000010111100:	sigmoid = 21'b000000000001111110111;
		14'b11000010111101:	sigmoid = 21'b000000000001111111001;
		14'b11000010111110:	sigmoid = 21'b000000000001111111011;
		14'b11000010111111:	sigmoid = 21'b000000000001111111101;
		14'b11000011000000:	sigmoid = 21'b000000000001111111111;
		14'b11000011000001:	sigmoid = 21'b000000000010000000001;
		14'b11000011000010:	sigmoid = 21'b000000000010000000011;
		14'b11000011000011:	sigmoid = 21'b000000000010000000101;
		14'b11000011000100:	sigmoid = 21'b000000000010000000111;
		14'b11000011000101:	sigmoid = 21'b000000000010000001001;
		14'b11000011000110:	sigmoid = 21'b000000000010000001011;
		14'b11000011000111:	sigmoid = 21'b000000000010000001101;
		14'b11000011001000:	sigmoid = 21'b000000000010000001111;
		14'b11000011001001:	sigmoid = 21'b000000000010000010001;
		14'b11000011001010:	sigmoid = 21'b000000000010000010011;
		14'b11000011001011:	sigmoid = 21'b000000000010000010101;
		14'b11000011001100:	sigmoid = 21'b000000000010000010111;
		14'b11000011001101:	sigmoid = 21'b000000000010000011001;
		14'b11000011001110:	sigmoid = 21'b000000000010000011011;
		14'b11000011001111:	sigmoid = 21'b000000000010000011101;
		14'b11000011010000:	sigmoid = 21'b000000000010000011111;
		14'b11000011010001:	sigmoid = 21'b000000000010000100001;
		14'b11000011010010:	sigmoid = 21'b000000000010000100011;
		14'b11000011010011:	sigmoid = 21'b000000000010000100101;
		14'b11000011010100:	sigmoid = 21'b000000000010000100111;
		14'b11000011010101:	sigmoid = 21'b000000000010000101001;
		14'b11000011010110:	sigmoid = 21'b000000000010000101100;
		14'b11000011010111:	sigmoid = 21'b000000000010000101110;
		14'b11000011011000:	sigmoid = 21'b000000000010000110000;
		14'b11000011011001:	sigmoid = 21'b000000000010000110010;
		14'b11000011011010:	sigmoid = 21'b000000000010000110100;
		14'b11000011011011:	sigmoid = 21'b000000000010000110110;
		14'b11000011011100:	sigmoid = 21'b000000000010000111000;
		14'b11000011011101:	sigmoid = 21'b000000000010000111010;
		14'b11000011011110:	sigmoid = 21'b000000000010000111100;
		14'b11000011011111:	sigmoid = 21'b000000000010000111110;
		14'b11000011100000:	sigmoid = 21'b000000000010001000001;
		14'b11000011100001:	sigmoid = 21'b000000000010001000011;
		14'b11000011100010:	sigmoid = 21'b000000000010001000101;
		14'b11000011100011:	sigmoid = 21'b000000000010001000111;
		14'b11000011100100:	sigmoid = 21'b000000000010001001001;
		14'b11000011100101:	sigmoid = 21'b000000000010001001011;
		14'b11000011100110:	sigmoid = 21'b000000000010001001101;
		14'b11000011100111:	sigmoid = 21'b000000000010001010000;
		14'b11000011101000:	sigmoid = 21'b000000000010001010010;
		14'b11000011101001:	sigmoid = 21'b000000000010001010100;
		14'b11000011101010:	sigmoid = 21'b000000000010001010110;
		14'b11000011101011:	sigmoid = 21'b000000000010001011000;
		14'b11000011101100:	sigmoid = 21'b000000000010001011010;
		14'b11000011101101:	sigmoid = 21'b000000000010001011101;
		14'b11000011101110:	sigmoid = 21'b000000000010001011111;
		14'b11000011101111:	sigmoid = 21'b000000000010001100001;
		14'b11000011110000:	sigmoid = 21'b000000000010001100011;
		14'b11000011110001:	sigmoid = 21'b000000000010001100101;
		14'b11000011110010:	sigmoid = 21'b000000000010001101000;
		14'b11000011110011:	sigmoid = 21'b000000000010001101010;
		14'b11000011110100:	sigmoid = 21'b000000000010001101100;
		14'b11000011110101:	sigmoid = 21'b000000000010001101110;
		14'b11000011110110:	sigmoid = 21'b000000000010001110000;
		14'b11000011110111:	sigmoid = 21'b000000000010001110011;
		14'b11000011111000:	sigmoid = 21'b000000000010001110101;
		14'b11000011111001:	sigmoid = 21'b000000000010001110111;
		14'b11000011111010:	sigmoid = 21'b000000000010001111001;
		14'b11000011111011:	sigmoid = 21'b000000000010001111100;
		14'b11000011111100:	sigmoid = 21'b000000000010001111110;
		14'b11000011111101:	sigmoid = 21'b000000000010010000000;
		14'b11000011111110:	sigmoid = 21'b000000000010010000010;
		14'b11000011111111:	sigmoid = 21'b000000000010010000101;
		14'b11000100000000:	sigmoid = 21'b000000000010010000111;
		14'b11000100000001:	sigmoid = 21'b000000000010010001001;
		14'b11000100000010:	sigmoid = 21'b000000000010010001011;
		14'b11000100000011:	sigmoid = 21'b000000000010010001110;
		14'b11000100000100:	sigmoid = 21'b000000000010010010000;
		14'b11000100000101:	sigmoid = 21'b000000000010010010010;
		14'b11000100000110:	sigmoid = 21'b000000000010010010100;
		14'b11000100000111:	sigmoid = 21'b000000000010010010111;
		14'b11000100001000:	sigmoid = 21'b000000000010010011001;
		14'b11000100001001:	sigmoid = 21'b000000000010010011011;
		14'b11000100001010:	sigmoid = 21'b000000000010010011110;
		14'b11000100001011:	sigmoid = 21'b000000000010010100000;
		14'b11000100001100:	sigmoid = 21'b000000000010010100010;
		14'b11000100001101:	sigmoid = 21'b000000000010010100101;
		14'b11000100001110:	sigmoid = 21'b000000000010010100111;
		14'b11000100001111:	sigmoid = 21'b000000000010010101001;
		14'b11000100010000:	sigmoid = 21'b000000000010010101100;
		14'b11000100010001:	sigmoid = 21'b000000000010010101110;
		14'b11000100010010:	sigmoid = 21'b000000000010010110000;
		14'b11000100010011:	sigmoid = 21'b000000000010010110011;
		14'b11000100010100:	sigmoid = 21'b000000000010010110101;
		14'b11000100010101:	sigmoid = 21'b000000000010010110111;
		14'b11000100010110:	sigmoid = 21'b000000000010010111010;
		14'b11000100010111:	sigmoid = 21'b000000000010010111100;
		14'b11000100011000:	sigmoid = 21'b000000000010010111110;
		14'b11000100011001:	sigmoid = 21'b000000000010011000001;
		14'b11000100011010:	sigmoid = 21'b000000000010011000011;
		14'b11000100011011:	sigmoid = 21'b000000000010011000101;
		14'b11000100011100:	sigmoid = 21'b000000000010011001000;
		14'b11000100011101:	sigmoid = 21'b000000000010011001010;
		14'b11000100011110:	sigmoid = 21'b000000000010011001101;
		14'b11000100011111:	sigmoid = 21'b000000000010011001111;
		14'b11000100100000:	sigmoid = 21'b000000000010011010001;
		14'b11000100100001:	sigmoid = 21'b000000000010011010100;
		14'b11000100100010:	sigmoid = 21'b000000000010011010110;
		14'b11000100100011:	sigmoid = 21'b000000000010011011001;
		14'b11000100100100:	sigmoid = 21'b000000000010011011011;
		14'b11000100100101:	sigmoid = 21'b000000000010011011110;
		14'b11000100100110:	sigmoid = 21'b000000000010011100000;
		14'b11000100100111:	sigmoid = 21'b000000000010011100010;
		14'b11000100101000:	sigmoid = 21'b000000000010011100101;
		14'b11000100101001:	sigmoid = 21'b000000000010011100111;
		14'b11000100101010:	sigmoid = 21'b000000000010011101010;
		14'b11000100101011:	sigmoid = 21'b000000000010011101100;
		14'b11000100101100:	sigmoid = 21'b000000000010011101111;
		14'b11000100101101:	sigmoid = 21'b000000000010011110001;
		14'b11000100101110:	sigmoid = 21'b000000000010011110100;
		14'b11000100101111:	sigmoid = 21'b000000000010011110110;
		14'b11000100110000:	sigmoid = 21'b000000000010011111001;
		14'b11000100110001:	sigmoid = 21'b000000000010011111011;
		14'b11000100110010:	sigmoid = 21'b000000000010011111110;
		14'b11000100110011:	sigmoid = 21'b000000000010100000000;
		14'b11000100110100:	sigmoid = 21'b000000000010100000011;
		14'b11000100110101:	sigmoid = 21'b000000000010100000101;
		14'b11000100110110:	sigmoid = 21'b000000000010100001000;
		14'b11000100110111:	sigmoid = 21'b000000000010100001010;
		14'b11000100111000:	sigmoid = 21'b000000000010100001101;
		14'b11000100111001:	sigmoid = 21'b000000000010100001111;
		14'b11000100111010:	sigmoid = 21'b000000000010100010010;
		14'b11000100111011:	sigmoid = 21'b000000000010100010100;
		14'b11000100111100:	sigmoid = 21'b000000000010100010111;
		14'b11000100111101:	sigmoid = 21'b000000000010100011001;
		14'b11000100111110:	sigmoid = 21'b000000000010100011100;
		14'b11000100111111:	sigmoid = 21'b000000000010100011110;
		14'b11000101000000:	sigmoid = 21'b000000000010100100001;
		14'b11000101000001:	sigmoid = 21'b000000000010100100100;
		14'b11000101000010:	sigmoid = 21'b000000000010100100110;
		14'b11000101000011:	sigmoid = 21'b000000000010100101001;
		14'b11000101000100:	sigmoid = 21'b000000000010100101011;
		14'b11000101000101:	sigmoid = 21'b000000000010100101110;
		14'b11000101000110:	sigmoid = 21'b000000000010100110000;
		14'b11000101000111:	sigmoid = 21'b000000000010100110011;
		14'b11000101001000:	sigmoid = 21'b000000000010100110110;
		14'b11000101001001:	sigmoid = 21'b000000000010100111000;
		14'b11000101001010:	sigmoid = 21'b000000000010100111011;
		14'b11000101001011:	sigmoid = 21'b000000000010100111110;
		14'b11000101001100:	sigmoid = 21'b000000000010101000000;
		14'b11000101001101:	sigmoid = 21'b000000000010101000011;
		14'b11000101001110:	sigmoid = 21'b000000000010101000101;
		14'b11000101001111:	sigmoid = 21'b000000000010101001000;
		14'b11000101010000:	sigmoid = 21'b000000000010101001011;
		14'b11000101010001:	sigmoid = 21'b000000000010101001101;
		14'b11000101010010:	sigmoid = 21'b000000000010101010000;
		14'b11000101010011:	sigmoid = 21'b000000000010101010011;
		14'b11000101010100:	sigmoid = 21'b000000000010101010101;
		14'b11000101010101:	sigmoid = 21'b000000000010101011000;
		14'b11000101010110:	sigmoid = 21'b000000000010101011011;
		14'b11000101010111:	sigmoid = 21'b000000000010101011101;
		14'b11000101011000:	sigmoid = 21'b000000000010101100000;
		14'b11000101011001:	sigmoid = 21'b000000000010101100011;
		14'b11000101011010:	sigmoid = 21'b000000000010101100101;
		14'b11000101011011:	sigmoid = 21'b000000000010101101000;
		14'b11000101011100:	sigmoid = 21'b000000000010101101011;
		14'b11000101011101:	sigmoid = 21'b000000000010101101110;
		14'b11000101011110:	sigmoid = 21'b000000000010101110000;
		14'b11000101011111:	sigmoid = 21'b000000000010101110011;
		14'b11000101100000:	sigmoid = 21'b000000000010101110110;
		14'b11000101100001:	sigmoid = 21'b000000000010101111000;
		14'b11000101100010:	sigmoid = 21'b000000000010101111011;
		14'b11000101100011:	sigmoid = 21'b000000000010101111110;
		14'b11000101100100:	sigmoid = 21'b000000000010110000001;
		14'b11000101100101:	sigmoid = 21'b000000000010110000011;
		14'b11000101100110:	sigmoid = 21'b000000000010110000110;
		14'b11000101100111:	sigmoid = 21'b000000000010110001001;
		14'b11000101101000:	sigmoid = 21'b000000000010110001100;
		14'b11000101101001:	sigmoid = 21'b000000000010110001110;
		14'b11000101101010:	sigmoid = 21'b000000000010110010001;
		14'b11000101101011:	sigmoid = 21'b000000000010110010100;
		14'b11000101101100:	sigmoid = 21'b000000000010110010111;
		14'b11000101101101:	sigmoid = 21'b000000000010110011010;
		14'b11000101101110:	sigmoid = 21'b000000000010110011100;
		14'b11000101101111:	sigmoid = 21'b000000000010110011111;
		14'b11000101110000:	sigmoid = 21'b000000000010110100010;
		14'b11000101110001:	sigmoid = 21'b000000000010110100101;
		14'b11000101110010:	sigmoid = 21'b000000000010110101000;
		14'b11000101110011:	sigmoid = 21'b000000000010110101010;
		14'b11000101110100:	sigmoid = 21'b000000000010110101101;
		14'b11000101110101:	sigmoid = 21'b000000000010110110000;
		14'b11000101110110:	sigmoid = 21'b000000000010110110011;
		14'b11000101110111:	sigmoid = 21'b000000000010110110110;
		14'b11000101111000:	sigmoid = 21'b000000000010110111001;
		14'b11000101111001:	sigmoid = 21'b000000000010110111100;
		14'b11000101111010:	sigmoid = 21'b000000000010110111110;
		14'b11000101111011:	sigmoid = 21'b000000000010111000001;
		14'b11000101111100:	sigmoid = 21'b000000000010111000100;
		14'b11000101111101:	sigmoid = 21'b000000000010111000111;
		14'b11000101111110:	sigmoid = 21'b000000000010111001010;
		14'b11000101111111:	sigmoid = 21'b000000000010111001101;
		14'b11000110000000:	sigmoid = 21'b000000000010111010000;
		14'b11000110000001:	sigmoid = 21'b000000000010111010011;
		14'b11000110000010:	sigmoid = 21'b000000000010111010110;
		14'b11000110000011:	sigmoid = 21'b000000000010111011001;
		14'b11000110000100:	sigmoid = 21'b000000000010111011011;
		14'b11000110000101:	sigmoid = 21'b000000000010111011110;
		14'b11000110000110:	sigmoid = 21'b000000000010111100001;
		14'b11000110000111:	sigmoid = 21'b000000000010111100100;
		14'b11000110001000:	sigmoid = 21'b000000000010111100111;
		14'b11000110001001:	sigmoid = 21'b000000000010111101010;
		14'b11000110001010:	sigmoid = 21'b000000000010111101101;
		14'b11000110001011:	sigmoid = 21'b000000000010111110000;
		14'b11000110001100:	sigmoid = 21'b000000000010111110011;
		14'b11000110001101:	sigmoid = 21'b000000000010111110110;
		14'b11000110001110:	sigmoid = 21'b000000000010111111001;
		14'b11000110001111:	sigmoid = 21'b000000000010111111100;
		14'b11000110010000:	sigmoid = 21'b000000000010111111111;
		14'b11000110010001:	sigmoid = 21'b000000000011000000010;
		14'b11000110010010:	sigmoid = 21'b000000000011000000101;
		14'b11000110010011:	sigmoid = 21'b000000000011000001000;
		14'b11000110010100:	sigmoid = 21'b000000000011000001011;
		14'b11000110010101:	sigmoid = 21'b000000000011000001110;
		14'b11000110010110:	sigmoid = 21'b000000000011000010001;
		14'b11000110010111:	sigmoid = 21'b000000000011000010100;
		14'b11000110011000:	sigmoid = 21'b000000000011000010111;
		14'b11000110011001:	sigmoid = 21'b000000000011000011010;
		14'b11000110011010:	sigmoid = 21'b000000000011000011101;
		14'b11000110011011:	sigmoid = 21'b000000000011000100000;
		14'b11000110011100:	sigmoid = 21'b000000000011000100011;
		14'b11000110011101:	sigmoid = 21'b000000000011000100110;
		14'b11000110011110:	sigmoid = 21'b000000000011000101010;
		14'b11000110011111:	sigmoid = 21'b000000000011000101101;
		14'b11000110100000:	sigmoid = 21'b000000000011000110000;
		14'b11000110100001:	sigmoid = 21'b000000000011000110011;
		14'b11000110100010:	sigmoid = 21'b000000000011000110110;
		14'b11000110100011:	sigmoid = 21'b000000000011000111001;
		14'b11000110100100:	sigmoid = 21'b000000000011000111100;
		14'b11000110100101:	sigmoid = 21'b000000000011000111111;
		14'b11000110100110:	sigmoid = 21'b000000000011001000010;
		14'b11000110100111:	sigmoid = 21'b000000000011001000101;
		14'b11000110101000:	sigmoid = 21'b000000000011001001001;
		14'b11000110101001:	sigmoid = 21'b000000000011001001100;
		14'b11000110101010:	sigmoid = 21'b000000000011001001111;
		14'b11000110101011:	sigmoid = 21'b000000000011001010010;
		14'b11000110101100:	sigmoid = 21'b000000000011001010101;
		14'b11000110101101:	sigmoid = 21'b000000000011001011000;
		14'b11000110101110:	sigmoid = 21'b000000000011001011100;
		14'b11000110101111:	sigmoid = 21'b000000000011001011111;
		14'b11000110110000:	sigmoid = 21'b000000000011001100010;
		14'b11000110110001:	sigmoid = 21'b000000000011001100101;
		14'b11000110110010:	sigmoid = 21'b000000000011001101000;
		14'b11000110110011:	sigmoid = 21'b000000000011001101100;
		14'b11000110110100:	sigmoid = 21'b000000000011001101111;
		14'b11000110110101:	sigmoid = 21'b000000000011001110010;
		14'b11000110110110:	sigmoid = 21'b000000000011001110101;
		14'b11000110110111:	sigmoid = 21'b000000000011001111000;
		14'b11000110111000:	sigmoid = 21'b000000000011001111100;
		14'b11000110111001:	sigmoid = 21'b000000000011001111111;
		14'b11000110111010:	sigmoid = 21'b000000000011010000010;
		14'b11000110111011:	sigmoid = 21'b000000000011010000101;
		14'b11000110111100:	sigmoid = 21'b000000000011010001001;
		14'b11000110111101:	sigmoid = 21'b000000000011010001100;
		14'b11000110111110:	sigmoid = 21'b000000000011010001111;
		14'b11000110111111:	sigmoid = 21'b000000000011010010011;
		14'b11000111000000:	sigmoid = 21'b000000000011010010110;
		14'b11000111000001:	sigmoid = 21'b000000000011010011001;
		14'b11000111000010:	sigmoid = 21'b000000000011010011100;
		14'b11000111000011:	sigmoid = 21'b000000000011010100000;
		14'b11000111000100:	sigmoid = 21'b000000000011010100011;
		14'b11000111000101:	sigmoid = 21'b000000000011010100110;
		14'b11000111000110:	sigmoid = 21'b000000000011010101010;
		14'b11000111000111:	sigmoid = 21'b000000000011010101101;
		14'b11000111001000:	sigmoid = 21'b000000000011010110000;
		14'b11000111001001:	sigmoid = 21'b000000000011010110100;
		14'b11000111001010:	sigmoid = 21'b000000000011010110111;
		14'b11000111001011:	sigmoid = 21'b000000000011010111010;
		14'b11000111001100:	sigmoid = 21'b000000000011010111110;
		14'b11000111001101:	sigmoid = 21'b000000000011011000001;
		14'b11000111001110:	sigmoid = 21'b000000000011011000100;
		14'b11000111001111:	sigmoid = 21'b000000000011011001000;
		14'b11000111010000:	sigmoid = 21'b000000000011011001011;
		14'b11000111010001:	sigmoid = 21'b000000000011011001111;
		14'b11000111010010:	sigmoid = 21'b000000000011011010010;
		14'b11000111010011:	sigmoid = 21'b000000000011011010101;
		14'b11000111010100:	sigmoid = 21'b000000000011011011001;
		14'b11000111010101:	sigmoid = 21'b000000000011011011100;
		14'b11000111010110:	sigmoid = 21'b000000000011011100000;
		14'b11000111010111:	sigmoid = 21'b000000000011011100011;
		14'b11000111011000:	sigmoid = 21'b000000000011011100111;
		14'b11000111011001:	sigmoid = 21'b000000000011011101010;
		14'b11000111011010:	sigmoid = 21'b000000000011011101110;
		14'b11000111011011:	sigmoid = 21'b000000000011011110001;
		14'b11000111011100:	sigmoid = 21'b000000000011011110100;
		14'b11000111011101:	sigmoid = 21'b000000000011011111000;
		14'b11000111011110:	sigmoid = 21'b000000000011011111011;
		14'b11000111011111:	sigmoid = 21'b000000000011011111111;
		14'b11000111100000:	sigmoid = 21'b000000000011100000010;
		14'b11000111100001:	sigmoid = 21'b000000000011100000110;
		14'b11000111100010:	sigmoid = 21'b000000000011100001001;
		14'b11000111100011:	sigmoid = 21'b000000000011100001101;
		14'b11000111100100:	sigmoid = 21'b000000000011100010001;
		14'b11000111100101:	sigmoid = 21'b000000000011100010100;
		14'b11000111100110:	sigmoid = 21'b000000000011100011000;
		14'b11000111100111:	sigmoid = 21'b000000000011100011011;
		14'b11000111101000:	sigmoid = 21'b000000000011100011111;
		14'b11000111101001:	sigmoid = 21'b000000000011100100010;
		14'b11000111101010:	sigmoid = 21'b000000000011100100110;
		14'b11000111101011:	sigmoid = 21'b000000000011100101001;
		14'b11000111101100:	sigmoid = 21'b000000000011100101101;
		14'b11000111101101:	sigmoid = 21'b000000000011100110001;
		14'b11000111101110:	sigmoid = 21'b000000000011100110100;
		14'b11000111101111:	sigmoid = 21'b000000000011100111000;
		14'b11000111110000:	sigmoid = 21'b000000000011100111011;
		14'b11000111110001:	sigmoid = 21'b000000000011100111111;
		14'b11000111110010:	sigmoid = 21'b000000000011101000011;
		14'b11000111110011:	sigmoid = 21'b000000000011101000110;
		14'b11000111110100:	sigmoid = 21'b000000000011101001010;
		14'b11000111110101:	sigmoid = 21'b000000000011101001110;
		14'b11000111110110:	sigmoid = 21'b000000000011101010001;
		14'b11000111110111:	sigmoid = 21'b000000000011101010101;
		14'b11000111111000:	sigmoid = 21'b000000000011101011001;
		14'b11000111111001:	sigmoid = 21'b000000000011101011100;
		14'b11000111111010:	sigmoid = 21'b000000000011101100000;
		14'b11000111111011:	sigmoid = 21'b000000000011101100100;
		14'b11000111111100:	sigmoid = 21'b000000000011101100111;
		14'b11000111111101:	sigmoid = 21'b000000000011101101011;
		14'b11000111111110:	sigmoid = 21'b000000000011101101111;
		14'b11000111111111:	sigmoid = 21'b000000000011101110010;
		14'b11001000000000:	sigmoid = 21'b000000000011101110110;
		14'b11001000000001:	sigmoid = 21'b000000000011101111010;
		14'b11001000000010:	sigmoid = 21'b000000000011101111110;
		14'b11001000000011:	sigmoid = 21'b000000000011110000001;
		14'b11001000000100:	sigmoid = 21'b000000000011110000101;
		14'b11001000000101:	sigmoid = 21'b000000000011110001001;
		14'b11001000000110:	sigmoid = 21'b000000000011110001101;
		14'b11001000000111:	sigmoid = 21'b000000000011110010000;
		14'b11001000001000:	sigmoid = 21'b000000000011110010100;
		14'b11001000001001:	sigmoid = 21'b000000000011110011000;
		14'b11001000001010:	sigmoid = 21'b000000000011110011100;
		14'b11001000001011:	sigmoid = 21'b000000000011110100000;
		14'b11001000001100:	sigmoid = 21'b000000000011110100011;
		14'b11001000001101:	sigmoid = 21'b000000000011110100111;
		14'b11001000001110:	sigmoid = 21'b000000000011110101011;
		14'b11001000001111:	sigmoid = 21'b000000000011110101111;
		14'b11001000010000:	sigmoid = 21'b000000000011110110011;
		14'b11001000010001:	sigmoid = 21'b000000000011110110111;
		14'b11001000010010:	sigmoid = 21'b000000000011110111010;
		14'b11001000010011:	sigmoid = 21'b000000000011110111110;
		14'b11001000010100:	sigmoid = 21'b000000000011111000010;
		14'b11001000010101:	sigmoid = 21'b000000000011111000110;
		14'b11001000010110:	sigmoid = 21'b000000000011111001010;
		14'b11001000010111:	sigmoid = 21'b000000000011111001110;
		14'b11001000011000:	sigmoid = 21'b000000000011111010010;
		14'b11001000011001:	sigmoid = 21'b000000000011111010110;
		14'b11001000011010:	sigmoid = 21'b000000000011111011010;
		14'b11001000011011:	sigmoid = 21'b000000000011111011101;
		14'b11001000011100:	sigmoid = 21'b000000000011111100001;
		14'b11001000011101:	sigmoid = 21'b000000000011111100101;
		14'b11001000011110:	sigmoid = 21'b000000000011111101001;
		14'b11001000011111:	sigmoid = 21'b000000000011111101101;
		14'b11001000100000:	sigmoid = 21'b000000000011111110001;
		14'b11001000100001:	sigmoid = 21'b000000000011111110101;
		14'b11001000100010:	sigmoid = 21'b000000000011111111001;
		14'b11001000100011:	sigmoid = 21'b000000000011111111101;
		14'b11001000100100:	sigmoid = 21'b000000000100000000001;
		14'b11001000100101:	sigmoid = 21'b000000000100000000101;
		14'b11001000100110:	sigmoid = 21'b000000000100000001001;
		14'b11001000100111:	sigmoid = 21'b000000000100000001101;
		14'b11001000101000:	sigmoid = 21'b000000000100000010001;
		14'b11001000101001:	sigmoid = 21'b000000000100000010101;
		14'b11001000101010:	sigmoid = 21'b000000000100000011001;
		14'b11001000101011:	sigmoid = 21'b000000000100000011101;
		14'b11001000101100:	sigmoid = 21'b000000000100000100001;
		14'b11001000101101:	sigmoid = 21'b000000000100000100101;
		14'b11001000101110:	sigmoid = 21'b000000000100000101010;
		14'b11001000101111:	sigmoid = 21'b000000000100000101110;
		14'b11001000110000:	sigmoid = 21'b000000000100000110010;
		14'b11001000110001:	sigmoid = 21'b000000000100000110110;
		14'b11001000110010:	sigmoid = 21'b000000000100000111010;
		14'b11001000110011:	sigmoid = 21'b000000000100000111110;
		14'b11001000110100:	sigmoid = 21'b000000000100001000010;
		14'b11001000110101:	sigmoid = 21'b000000000100001000110;
		14'b11001000110110:	sigmoid = 21'b000000000100001001010;
		14'b11001000110111:	sigmoid = 21'b000000000100001001111;
		14'b11001000111000:	sigmoid = 21'b000000000100001010011;
		14'b11001000111001:	sigmoid = 21'b000000000100001010111;
		14'b11001000111010:	sigmoid = 21'b000000000100001011011;
		14'b11001000111011:	sigmoid = 21'b000000000100001011111;
		14'b11001000111100:	sigmoid = 21'b000000000100001100011;
		14'b11001000111101:	sigmoid = 21'b000000000100001101000;
		14'b11001000111110:	sigmoid = 21'b000000000100001101100;
		14'b11001000111111:	sigmoid = 21'b000000000100001110000;
		14'b11001001000000:	sigmoid = 21'b000000000100001110100;
		14'b11001001000001:	sigmoid = 21'b000000000100001111000;
		14'b11001001000010:	sigmoid = 21'b000000000100001111101;
		14'b11001001000011:	sigmoid = 21'b000000000100010000001;
		14'b11001001000100:	sigmoid = 21'b000000000100010000101;
		14'b11001001000101:	sigmoid = 21'b000000000100010001001;
		14'b11001001000110:	sigmoid = 21'b000000000100010001110;
		14'b11001001000111:	sigmoid = 21'b000000000100010010010;
		14'b11001001001000:	sigmoid = 21'b000000000100010010110;
		14'b11001001001001:	sigmoid = 21'b000000000100010011011;
		14'b11001001001010:	sigmoid = 21'b000000000100010011111;
		14'b11001001001011:	sigmoid = 21'b000000000100010100011;
		14'b11001001001100:	sigmoid = 21'b000000000100010101000;
		14'b11001001001101:	sigmoid = 21'b000000000100010101100;
		14'b11001001001110:	sigmoid = 21'b000000000100010110000;
		14'b11001001001111:	sigmoid = 21'b000000000100010110101;
		14'b11001001010000:	sigmoid = 21'b000000000100010111001;
		14'b11001001010001:	sigmoid = 21'b000000000100010111101;
		14'b11001001010010:	sigmoid = 21'b000000000100011000010;
		14'b11001001010011:	sigmoid = 21'b000000000100011000110;
		14'b11001001010100:	sigmoid = 21'b000000000100011001010;
		14'b11001001010101:	sigmoid = 21'b000000000100011001111;
		14'b11001001010110:	sigmoid = 21'b000000000100011010011;
		14'b11001001010111:	sigmoid = 21'b000000000100011011000;
		14'b11001001011000:	sigmoid = 21'b000000000100011011100;
		14'b11001001011001:	sigmoid = 21'b000000000100011100000;
		14'b11001001011010:	sigmoid = 21'b000000000100011100101;
		14'b11001001011011:	sigmoid = 21'b000000000100011101001;
		14'b11001001011100:	sigmoid = 21'b000000000100011101110;
		14'b11001001011101:	sigmoid = 21'b000000000100011110010;
		14'b11001001011110:	sigmoid = 21'b000000000100011110111;
		14'b11001001011111:	sigmoid = 21'b000000000100011111011;
		14'b11001001100000:	sigmoid = 21'b000000000100100000000;
		14'b11001001100001:	sigmoid = 21'b000000000100100000100;
		14'b11001001100010:	sigmoid = 21'b000000000100100001001;
		14'b11001001100011:	sigmoid = 21'b000000000100100001101;
		14'b11001001100100:	sigmoid = 21'b000000000100100010010;
		14'b11001001100101:	sigmoid = 21'b000000000100100010110;
		14'b11001001100110:	sigmoid = 21'b000000000100100011011;
		14'b11001001100111:	sigmoid = 21'b000000000100100011111;
		14'b11001001101000:	sigmoid = 21'b000000000100100100100;
		14'b11001001101001:	sigmoid = 21'b000000000100100101001;
		14'b11001001101010:	sigmoid = 21'b000000000100100101101;
		14'b11001001101011:	sigmoid = 21'b000000000100100110010;
		14'b11001001101100:	sigmoid = 21'b000000000100100110110;
		14'b11001001101101:	sigmoid = 21'b000000000100100111011;
		14'b11001001101110:	sigmoid = 21'b000000000100101000000;
		14'b11001001101111:	sigmoid = 21'b000000000100101000100;
		14'b11001001110000:	sigmoid = 21'b000000000100101001001;
		14'b11001001110001:	sigmoid = 21'b000000000100101001101;
		14'b11001001110010:	sigmoid = 21'b000000000100101010010;
		14'b11001001110011:	sigmoid = 21'b000000000100101010111;
		14'b11001001110100:	sigmoid = 21'b000000000100101011011;
		14'b11001001110101:	sigmoid = 21'b000000000100101100000;
		14'b11001001110110:	sigmoid = 21'b000000000100101100101;
		14'b11001001110111:	sigmoid = 21'b000000000100101101001;
		14'b11001001111000:	sigmoid = 21'b000000000100101101110;
		14'b11001001111001:	sigmoid = 21'b000000000100101110011;
		14'b11001001111010:	sigmoid = 21'b000000000100101111000;
		14'b11001001111011:	sigmoid = 21'b000000000100101111100;
		14'b11001001111100:	sigmoid = 21'b000000000100110000001;
		14'b11001001111101:	sigmoid = 21'b000000000100110000110;
		14'b11001001111110:	sigmoid = 21'b000000000100110001011;
		14'b11001001111111:	sigmoid = 21'b000000000100110001111;
		14'b11001010000000:	sigmoid = 21'b000000000100110010100;
		14'b11001010000001:	sigmoid = 21'b000000000100110011001;
		14'b11001010000010:	sigmoid = 21'b000000000100110011110;
		14'b11001010000011:	sigmoid = 21'b000000000100110100011;
		14'b11001010000100:	sigmoid = 21'b000000000100110100111;
		14'b11001010000101:	sigmoid = 21'b000000000100110101100;
		14'b11001010000110:	sigmoid = 21'b000000000100110110001;
		14'b11001010000111:	sigmoid = 21'b000000000100110110110;
		14'b11001010001000:	sigmoid = 21'b000000000100110111011;
		14'b11001010001001:	sigmoid = 21'b000000000100111000000;
		14'b11001010001010:	sigmoid = 21'b000000000100111000100;
		14'b11001010001011:	sigmoid = 21'b000000000100111001001;
		14'b11001010001100:	sigmoid = 21'b000000000100111001110;
		14'b11001010001101:	sigmoid = 21'b000000000100111010011;
		14'b11001010001110:	sigmoid = 21'b000000000100111011000;
		14'b11001010001111:	sigmoid = 21'b000000000100111011101;
		14'b11001010010000:	sigmoid = 21'b000000000100111100010;
		14'b11001010010001:	sigmoid = 21'b000000000100111100111;
		14'b11001010010010:	sigmoid = 21'b000000000100111101100;
		14'b11001010010011:	sigmoid = 21'b000000000100111110001;
		14'b11001010010100:	sigmoid = 21'b000000000100111110110;
		14'b11001010010101:	sigmoid = 21'b000000000100111111011;
		14'b11001010010110:	sigmoid = 21'b000000000101000000000;
		14'b11001010010111:	sigmoid = 21'b000000000101000000101;
		14'b11001010011000:	sigmoid = 21'b000000000101000001010;
		14'b11001010011001:	sigmoid = 21'b000000000101000001111;
		14'b11001010011010:	sigmoid = 21'b000000000101000010100;
		14'b11001010011011:	sigmoid = 21'b000000000101000011001;
		14'b11001010011100:	sigmoid = 21'b000000000101000011110;
		14'b11001010011101:	sigmoid = 21'b000000000101000100011;
		14'b11001010011110:	sigmoid = 21'b000000000101000101000;
		14'b11001010011111:	sigmoid = 21'b000000000101000101101;
		14'b11001010100000:	sigmoid = 21'b000000000101000110010;
		14'b11001010100001:	sigmoid = 21'b000000000101000110111;
		14'b11001010100010:	sigmoid = 21'b000000000101000111100;
		14'b11001010100011:	sigmoid = 21'b000000000101001000001;
		14'b11001010100100:	sigmoid = 21'b000000000101001000111;
		14'b11001010100101:	sigmoid = 21'b000000000101001001100;
		14'b11001010100110:	sigmoid = 21'b000000000101001010001;
		14'b11001010100111:	sigmoid = 21'b000000000101001010110;
		14'b11001010101000:	sigmoid = 21'b000000000101001011011;
		14'b11001010101001:	sigmoid = 21'b000000000101001100000;
		14'b11001010101010:	sigmoid = 21'b000000000101001100110;
		14'b11001010101011:	sigmoid = 21'b000000000101001101011;
		14'b11001010101100:	sigmoid = 21'b000000000101001110000;
		14'b11001010101101:	sigmoid = 21'b000000000101001110101;
		14'b11001010101110:	sigmoid = 21'b000000000101001111010;
		14'b11001010101111:	sigmoid = 21'b000000000101010000000;
		14'b11001010110000:	sigmoid = 21'b000000000101010000101;
		14'b11001010110001:	sigmoid = 21'b000000000101010001010;
		14'b11001010110010:	sigmoid = 21'b000000000101010001111;
		14'b11001010110011:	sigmoid = 21'b000000000101010010101;
		14'b11001010110100:	sigmoid = 21'b000000000101010011010;
		14'b11001010110101:	sigmoid = 21'b000000000101010011111;
		14'b11001010110110:	sigmoid = 21'b000000000101010100101;
		14'b11001010110111:	sigmoid = 21'b000000000101010101010;
		14'b11001010111000:	sigmoid = 21'b000000000101010101111;
		14'b11001010111001:	sigmoid = 21'b000000000101010110101;
		14'b11001010111010:	sigmoid = 21'b000000000101010111010;
		14'b11001010111011:	sigmoid = 21'b000000000101010111111;
		14'b11001010111100:	sigmoid = 21'b000000000101011000101;
		14'b11001010111101:	sigmoid = 21'b000000000101011001010;
		14'b11001010111110:	sigmoid = 21'b000000000101011001111;
		14'b11001010111111:	sigmoid = 21'b000000000101011010101;
		14'b11001011000000:	sigmoid = 21'b000000000101011011010;
		14'b11001011000001:	sigmoid = 21'b000000000101011100000;
		14'b11001011000010:	sigmoid = 21'b000000000101011100101;
		14'b11001011000011:	sigmoid = 21'b000000000101011101011;
		14'b11001011000100:	sigmoid = 21'b000000000101011110000;
		14'b11001011000101:	sigmoid = 21'b000000000101011110110;
		14'b11001011000110:	sigmoid = 21'b000000000101011111011;
		14'b11001011000111:	sigmoid = 21'b000000000101100000000;
		14'b11001011001000:	sigmoid = 21'b000000000101100000110;
		14'b11001011001001:	sigmoid = 21'b000000000101100001011;
		14'b11001011001010:	sigmoid = 21'b000000000101100010001;
		14'b11001011001011:	sigmoid = 21'b000000000101100010111;
		14'b11001011001100:	sigmoid = 21'b000000000101100011100;
		14'b11001011001101:	sigmoid = 21'b000000000101100100010;
		14'b11001011001110:	sigmoid = 21'b000000000101100100111;
		14'b11001011001111:	sigmoid = 21'b000000000101100101101;
		14'b11001011010000:	sigmoid = 21'b000000000101100110010;
		14'b11001011010001:	sigmoid = 21'b000000000101100111000;
		14'b11001011010010:	sigmoid = 21'b000000000101100111110;
		14'b11001011010011:	sigmoid = 21'b000000000101101000011;
		14'b11001011010100:	sigmoid = 21'b000000000101101001001;
		14'b11001011010101:	sigmoid = 21'b000000000101101001110;
		14'b11001011010110:	sigmoid = 21'b000000000101101010100;
		14'b11001011010111:	sigmoid = 21'b000000000101101011010;
		14'b11001011011000:	sigmoid = 21'b000000000101101011111;
		14'b11001011011001:	sigmoid = 21'b000000000101101100101;
		14'b11001011011010:	sigmoid = 21'b000000000101101101011;
		14'b11001011011011:	sigmoid = 21'b000000000101101110001;
		14'b11001011011100:	sigmoid = 21'b000000000101101110110;
		14'b11001011011101:	sigmoid = 21'b000000000101101111100;
		14'b11001011011110:	sigmoid = 21'b000000000101110000010;
		14'b11001011011111:	sigmoid = 21'b000000000101110000111;
		14'b11001011100000:	sigmoid = 21'b000000000101110001101;
		14'b11001011100001:	sigmoid = 21'b000000000101110010011;
		14'b11001011100010:	sigmoid = 21'b000000000101110011001;
		14'b11001011100011:	sigmoid = 21'b000000000101110011111;
		14'b11001011100100:	sigmoid = 21'b000000000101110100100;
		14'b11001011100101:	sigmoid = 21'b000000000101110101010;
		14'b11001011100110:	sigmoid = 21'b000000000101110110000;
		14'b11001011100111:	sigmoid = 21'b000000000101110110110;
		14'b11001011101000:	sigmoid = 21'b000000000101110111100;
		14'b11001011101001:	sigmoid = 21'b000000000101111000010;
		14'b11001011101010:	sigmoid = 21'b000000000101111000111;
		14'b11001011101011:	sigmoid = 21'b000000000101111001101;
		14'b11001011101100:	sigmoid = 21'b000000000101111010011;
		14'b11001011101101:	sigmoid = 21'b000000000101111011001;
		14'b11001011101110:	sigmoid = 21'b000000000101111011111;
		14'b11001011101111:	sigmoid = 21'b000000000101111100101;
		14'b11001011110000:	sigmoid = 21'b000000000101111101011;
		14'b11001011110001:	sigmoid = 21'b000000000101111110001;
		14'b11001011110010:	sigmoid = 21'b000000000101111110111;
		14'b11001011110011:	sigmoid = 21'b000000000101111111101;
		14'b11001011110100:	sigmoid = 21'b000000000110000000011;
		14'b11001011110101:	sigmoid = 21'b000000000110000001001;
		14'b11001011110110:	sigmoid = 21'b000000000110000001111;
		14'b11001011110111:	sigmoid = 21'b000000000110000010101;
		14'b11001011111000:	sigmoid = 21'b000000000110000011011;
		14'b11001011111001:	sigmoid = 21'b000000000110000100001;
		14'b11001011111010:	sigmoid = 21'b000000000110000100111;
		14'b11001011111011:	sigmoid = 21'b000000000110000101101;
		14'b11001011111100:	sigmoid = 21'b000000000110000110011;
		14'b11001011111101:	sigmoid = 21'b000000000110000111001;
		14'b11001011111110:	sigmoid = 21'b000000000110000111111;
		14'b11001011111111:	sigmoid = 21'b000000000110001000110;
		14'b11001100000000:	sigmoid = 21'b000000000110001001100;
		14'b11001100000001:	sigmoid = 21'b000000000110001010010;
		14'b11001100000010:	sigmoid = 21'b000000000110001011000;
		14'b11001100000011:	sigmoid = 21'b000000000110001011110;
		14'b11001100000100:	sigmoid = 21'b000000000110001100100;
		14'b11001100000101:	sigmoid = 21'b000000000110001101011;
		14'b11001100000110:	sigmoid = 21'b000000000110001110001;
		14'b11001100000111:	sigmoid = 21'b000000000110001110111;
		14'b11001100001000:	sigmoid = 21'b000000000110001111101;
		14'b11001100001001:	sigmoid = 21'b000000000110010000011;
		14'b11001100001010:	sigmoid = 21'b000000000110010001010;
		14'b11001100001011:	sigmoid = 21'b000000000110010010000;
		14'b11001100001100:	sigmoid = 21'b000000000110010010110;
		14'b11001100001101:	sigmoid = 21'b000000000110010011101;
		14'b11001100001110:	sigmoid = 21'b000000000110010100011;
		14'b11001100001111:	sigmoid = 21'b000000000110010101001;
		14'b11001100010000:	sigmoid = 21'b000000000110010101111;
		14'b11001100010001:	sigmoid = 21'b000000000110010110110;
		14'b11001100010010:	sigmoid = 21'b000000000110010111100;
		14'b11001100010011:	sigmoid = 21'b000000000110011000011;
		14'b11001100010100:	sigmoid = 21'b000000000110011001001;
		14'b11001100010101:	sigmoid = 21'b000000000110011001111;
		14'b11001100010110:	sigmoid = 21'b000000000110011010110;
		14'b11001100010111:	sigmoid = 21'b000000000110011011100;
		14'b11001100011000:	sigmoid = 21'b000000000110011100011;
		14'b11001100011001:	sigmoid = 21'b000000000110011101001;
		14'b11001100011010:	sigmoid = 21'b000000000110011101111;
		14'b11001100011011:	sigmoid = 21'b000000000110011110110;
		14'b11001100011100:	sigmoid = 21'b000000000110011111100;
		14'b11001100011101:	sigmoid = 21'b000000000110100000011;
		14'b11001100011110:	sigmoid = 21'b000000000110100001001;
		14'b11001100011111:	sigmoid = 21'b000000000110100010000;
		14'b11001100100000:	sigmoid = 21'b000000000110100010110;
		14'b11001100100001:	sigmoid = 21'b000000000110100011101;
		14'b11001100100010:	sigmoid = 21'b000000000110100100100;
		14'b11001100100011:	sigmoid = 21'b000000000110100101010;
		14'b11001100100100:	sigmoid = 21'b000000000110100110001;
		14'b11001100100101:	sigmoid = 21'b000000000110100110111;
		14'b11001100100110:	sigmoid = 21'b000000000110100111110;
		14'b11001100100111:	sigmoid = 21'b000000000110101000100;
		14'b11001100101000:	sigmoid = 21'b000000000110101001011;
		14'b11001100101001:	sigmoid = 21'b000000000110101010010;
		14'b11001100101010:	sigmoid = 21'b000000000110101011000;
		14'b11001100101011:	sigmoid = 21'b000000000110101011111;
		14'b11001100101100:	sigmoid = 21'b000000000110101100110;
		14'b11001100101101:	sigmoid = 21'b000000000110101101100;
		14'b11001100101110:	sigmoid = 21'b000000000110101110011;
		14'b11001100101111:	sigmoid = 21'b000000000110101111010;
		14'b11001100110000:	sigmoid = 21'b000000000110110000001;
		14'b11001100110001:	sigmoid = 21'b000000000110110000111;
		14'b11001100110010:	sigmoid = 21'b000000000110110001110;
		14'b11001100110011:	sigmoid = 21'b000000000110110010101;
		14'b11001100110100:	sigmoid = 21'b000000000110110011100;
		14'b11001100110101:	sigmoid = 21'b000000000110110100010;
		14'b11001100110110:	sigmoid = 21'b000000000110110101001;
		14'b11001100110111:	sigmoid = 21'b000000000110110110000;
		14'b11001100111000:	sigmoid = 21'b000000000110110110111;
		14'b11001100111001:	sigmoid = 21'b000000000110110111110;
		14'b11001100111010:	sigmoid = 21'b000000000110111000101;
		14'b11001100111011:	sigmoid = 21'b000000000110111001100;
		14'b11001100111100:	sigmoid = 21'b000000000110111010010;
		14'b11001100111101:	sigmoid = 21'b000000000110111011001;
		14'b11001100111110:	sigmoid = 21'b000000000110111100000;
		14'b11001100111111:	sigmoid = 21'b000000000110111100111;
		14'b11001101000000:	sigmoid = 21'b000000000110111101110;
		14'b11001101000001:	sigmoid = 21'b000000000110111110101;
		14'b11001101000010:	sigmoid = 21'b000000000110111111100;
		14'b11001101000011:	sigmoid = 21'b000000000111000000011;
		14'b11001101000100:	sigmoid = 21'b000000000111000001010;
		14'b11001101000101:	sigmoid = 21'b000000000111000010001;
		14'b11001101000110:	sigmoid = 21'b000000000111000011000;
		14'b11001101000111:	sigmoid = 21'b000000000111000011111;
		14'b11001101001000:	sigmoid = 21'b000000000111000100110;
		14'b11001101001001:	sigmoid = 21'b000000000111000101101;
		14'b11001101001010:	sigmoid = 21'b000000000111000110100;
		14'b11001101001011:	sigmoid = 21'b000000000111000111011;
		14'b11001101001100:	sigmoid = 21'b000000000111001000011;
		14'b11001101001101:	sigmoid = 21'b000000000111001001010;
		14'b11001101001110:	sigmoid = 21'b000000000111001010001;
		14'b11001101001111:	sigmoid = 21'b000000000111001011000;
		14'b11001101010000:	sigmoid = 21'b000000000111001011111;
		14'b11001101010001:	sigmoid = 21'b000000000111001100110;
		14'b11001101010010:	sigmoid = 21'b000000000111001101110;
		14'b11001101010011:	sigmoid = 21'b000000000111001110101;
		14'b11001101010100:	sigmoid = 21'b000000000111001111100;
		14'b11001101010101:	sigmoid = 21'b000000000111010000011;
		14'b11001101010110:	sigmoid = 21'b000000000111010001010;
		14'b11001101010111:	sigmoid = 21'b000000000111010010010;
		14'b11001101011000:	sigmoid = 21'b000000000111010011001;
		14'b11001101011001:	sigmoid = 21'b000000000111010100000;
		14'b11001101011010:	sigmoid = 21'b000000000111010101000;
		14'b11001101011011:	sigmoid = 21'b000000000111010101111;
		14'b11001101011100:	sigmoid = 21'b000000000111010110110;
		14'b11001101011101:	sigmoid = 21'b000000000111010111110;
		14'b11001101011110:	sigmoid = 21'b000000000111011000101;
		14'b11001101011111:	sigmoid = 21'b000000000111011001100;
		14'b11001101100000:	sigmoid = 21'b000000000111011010100;
		14'b11001101100001:	sigmoid = 21'b000000000111011011011;
		14'b11001101100010:	sigmoid = 21'b000000000111011100011;
		14'b11001101100011:	sigmoid = 21'b000000000111011101010;
		14'b11001101100100:	sigmoid = 21'b000000000111011110010;
		14'b11001101100101:	sigmoid = 21'b000000000111011111001;
		14'b11001101100110:	sigmoid = 21'b000000000111100000000;
		14'b11001101100111:	sigmoid = 21'b000000000111100001000;
		14'b11001101101000:	sigmoid = 21'b000000000111100001111;
		14'b11001101101001:	sigmoid = 21'b000000000111100010111;
		14'b11001101101010:	sigmoid = 21'b000000000111100011111;
		14'b11001101101011:	sigmoid = 21'b000000000111100100110;
		14'b11001101101100:	sigmoid = 21'b000000000111100101110;
		14'b11001101101101:	sigmoid = 21'b000000000111100110101;
		14'b11001101101110:	sigmoid = 21'b000000000111100111101;
		14'b11001101101111:	sigmoid = 21'b000000000111101000100;
		14'b11001101110000:	sigmoid = 21'b000000000111101001100;
		14'b11001101110001:	sigmoid = 21'b000000000111101010100;
		14'b11001101110010:	sigmoid = 21'b000000000111101011011;
		14'b11001101110011:	sigmoid = 21'b000000000111101100011;
		14'b11001101110100:	sigmoid = 21'b000000000111101101011;
		14'b11001101110101:	sigmoid = 21'b000000000111101110010;
		14'b11001101110110:	sigmoid = 21'b000000000111101111010;
		14'b11001101110111:	sigmoid = 21'b000000000111110000010;
		14'b11001101111000:	sigmoid = 21'b000000000111110001010;
		14'b11001101111001:	sigmoid = 21'b000000000111110010001;
		14'b11001101111010:	sigmoid = 21'b000000000111110011001;
		14'b11001101111011:	sigmoid = 21'b000000000111110100001;
		14'b11001101111100:	sigmoid = 21'b000000000111110101001;
		14'b11001101111101:	sigmoid = 21'b000000000111110110001;
		14'b11001101111110:	sigmoid = 21'b000000000111110111000;
		14'b11001101111111:	sigmoid = 21'b000000000111111000000;
		14'b11001110000000:	sigmoid = 21'b000000000111111001000;
		14'b11001110000001:	sigmoid = 21'b000000000111111010000;
		14'b11001110000010:	sigmoid = 21'b000000000111111011000;
		14'b11001110000011:	sigmoid = 21'b000000000111111100000;
		14'b11001110000100:	sigmoid = 21'b000000000111111101000;
		14'b11001110000101:	sigmoid = 21'b000000000111111110000;
		14'b11001110000110:	sigmoid = 21'b000000000111111111000;
		14'b11001110000111:	sigmoid = 21'b000000001000000000000;
		14'b11001110001000:	sigmoid = 21'b000000001000000001000;
		14'b11001110001001:	sigmoid = 21'b000000001000000010000;
		14'b11001110001010:	sigmoid = 21'b000000001000000011000;
		14'b11001110001011:	sigmoid = 21'b000000001000000100000;
		14'b11001110001100:	sigmoid = 21'b000000001000000101000;
		14'b11001110001101:	sigmoid = 21'b000000001000000110000;
		14'b11001110001110:	sigmoid = 21'b000000001000000111000;
		14'b11001110001111:	sigmoid = 21'b000000001000001000000;
		14'b11001110010000:	sigmoid = 21'b000000001000001001000;
		14'b11001110010001:	sigmoid = 21'b000000001000001010000;
		14'b11001110010010:	sigmoid = 21'b000000001000001011000;
		14'b11001110010011:	sigmoid = 21'b000000001000001100001;
		14'b11001110010100:	sigmoid = 21'b000000001000001101001;
		14'b11001110010101:	sigmoid = 21'b000000001000001110001;
		14'b11001110010110:	sigmoid = 21'b000000001000001111001;
		14'b11001110010111:	sigmoid = 21'b000000001000010000001;
		14'b11001110011000:	sigmoid = 21'b000000001000010001010;
		14'b11001110011001:	sigmoid = 21'b000000001000010010010;
		14'b11001110011010:	sigmoid = 21'b000000001000010011010;
		14'b11001110011011:	sigmoid = 21'b000000001000010100011;
		14'b11001110011100:	sigmoid = 21'b000000001000010101011;
		14'b11001110011101:	sigmoid = 21'b000000001000010110011;
		14'b11001110011110:	sigmoid = 21'b000000001000010111011;
		14'b11001110011111:	sigmoid = 21'b000000001000011000100;
		14'b11001110100000:	sigmoid = 21'b000000001000011001100;
		14'b11001110100001:	sigmoid = 21'b000000001000011010101;
		14'b11001110100010:	sigmoid = 21'b000000001000011011101;
		14'b11001110100011:	sigmoid = 21'b000000001000011100101;
		14'b11001110100100:	sigmoid = 21'b000000001000011101110;
		14'b11001110100101:	sigmoid = 21'b000000001000011110110;
		14'b11001110100110:	sigmoid = 21'b000000001000011111111;
		14'b11001110100111:	sigmoid = 21'b000000001000100000111;
		14'b11001110101000:	sigmoid = 21'b000000001000100010000;
		14'b11001110101001:	sigmoid = 21'b000000001000100011000;
		14'b11001110101010:	sigmoid = 21'b000000001000100100001;
		14'b11001110101011:	sigmoid = 21'b000000001000100101001;
		14'b11001110101100:	sigmoid = 21'b000000001000100110010;
		14'b11001110101101:	sigmoid = 21'b000000001000100111011;
		14'b11001110101110:	sigmoid = 21'b000000001000101000011;
		14'b11001110101111:	sigmoid = 21'b000000001000101001100;
		14'b11001110110000:	sigmoid = 21'b000000001000101010100;
		14'b11001110110001:	sigmoid = 21'b000000001000101011101;
		14'b11001110110010:	sigmoid = 21'b000000001000101100110;
		14'b11001110110011:	sigmoid = 21'b000000001000101101110;
		14'b11001110110100:	sigmoid = 21'b000000001000101110111;
		14'b11001110110101:	sigmoid = 21'b000000001000110000000;
		14'b11001110110110:	sigmoid = 21'b000000001000110001001;
		14'b11001110110111:	sigmoid = 21'b000000001000110010001;
		14'b11001110111000:	sigmoid = 21'b000000001000110011010;
		14'b11001110111001:	sigmoid = 21'b000000001000110100011;
		14'b11001110111010:	sigmoid = 21'b000000001000110101100;
		14'b11001110111011:	sigmoid = 21'b000000001000110110101;
		14'b11001110111100:	sigmoid = 21'b000000001000110111101;
		14'b11001110111101:	sigmoid = 21'b000000001000111000110;
		14'b11001110111110:	sigmoid = 21'b000000001000111001111;
		14'b11001110111111:	sigmoid = 21'b000000001000111011000;
		14'b11001111000000:	sigmoid = 21'b000000001000111100001;
		14'b11001111000001:	sigmoid = 21'b000000001000111101010;
		14'b11001111000010:	sigmoid = 21'b000000001000111110011;
		14'b11001111000011:	sigmoid = 21'b000000001000111111100;
		14'b11001111000100:	sigmoid = 21'b000000001001000000101;
		14'b11001111000101:	sigmoid = 21'b000000001001000001110;
		14'b11001111000110:	sigmoid = 21'b000000001001000010111;
		14'b11001111000111:	sigmoid = 21'b000000001001000100000;
		14'b11001111001000:	sigmoid = 21'b000000001001000101001;
		14'b11001111001001:	sigmoid = 21'b000000001001000110010;
		14'b11001111001010:	sigmoid = 21'b000000001001000111011;
		14'b11001111001011:	sigmoid = 21'b000000001001001000100;
		14'b11001111001100:	sigmoid = 21'b000000001001001001101;
		14'b11001111001101:	sigmoid = 21'b000000001001001010110;
		14'b11001111001110:	sigmoid = 21'b000000001001001100000;
		14'b11001111001111:	sigmoid = 21'b000000001001001101001;
		14'b11001111010000:	sigmoid = 21'b000000001001001110010;
		14'b11001111010001:	sigmoid = 21'b000000001001001111011;
		14'b11001111010010:	sigmoid = 21'b000000001001010000100;
		14'b11001111010011:	sigmoid = 21'b000000001001010001110;
		14'b11001111010100:	sigmoid = 21'b000000001001010010111;
		14'b11001111010101:	sigmoid = 21'b000000001001010100000;
		14'b11001111010110:	sigmoid = 21'b000000001001010101010;
		14'b11001111010111:	sigmoid = 21'b000000001001010110011;
		14'b11001111011000:	sigmoid = 21'b000000001001010111100;
		14'b11001111011001:	sigmoid = 21'b000000001001011000110;
		14'b11001111011010:	sigmoid = 21'b000000001001011001111;
		14'b11001111011011:	sigmoid = 21'b000000001001011011000;
		14'b11001111011100:	sigmoid = 21'b000000001001011100010;
		14'b11001111011101:	sigmoid = 21'b000000001001011101011;
		14'b11001111011110:	sigmoid = 21'b000000001001011110101;
		14'b11001111011111:	sigmoid = 21'b000000001001011111110;
		14'b11001111100000:	sigmoid = 21'b000000001001100001000;
		14'b11001111100001:	sigmoid = 21'b000000001001100010001;
		14'b11001111100010:	sigmoid = 21'b000000001001100011011;
		14'b11001111100011:	sigmoid = 21'b000000001001100100100;
		14'b11001111100100:	sigmoid = 21'b000000001001100101110;
		14'b11001111100101:	sigmoid = 21'b000000001001100110111;
		14'b11001111100110:	sigmoid = 21'b000000001001101000001;
		14'b11001111100111:	sigmoid = 21'b000000001001101001010;
		14'b11001111101000:	sigmoid = 21'b000000001001101010100;
		14'b11001111101001:	sigmoid = 21'b000000001001101011110;
		14'b11001111101010:	sigmoid = 21'b000000001001101100111;
		14'b11001111101011:	sigmoid = 21'b000000001001101110001;
		14'b11001111101100:	sigmoid = 21'b000000001001101111011;
		14'b11001111101101:	sigmoid = 21'b000000001001110000101;
		14'b11001111101110:	sigmoid = 21'b000000001001110001110;
		14'b11001111101111:	sigmoid = 21'b000000001001110011000;
		14'b11001111110000:	sigmoid = 21'b000000001001110100010;
		14'b11001111110001:	sigmoid = 21'b000000001001110101100;
		14'b11001111110010:	sigmoid = 21'b000000001001110110101;
		14'b11001111110011:	sigmoid = 21'b000000001001110111111;
		14'b11001111110100:	sigmoid = 21'b000000001001111001001;
		14'b11001111110101:	sigmoid = 21'b000000001001111010011;
		14'b11001111110110:	sigmoid = 21'b000000001001111011101;
		14'b11001111110111:	sigmoid = 21'b000000001001111100111;
		14'b11001111111000:	sigmoid = 21'b000000001001111110001;
		14'b11001111111001:	sigmoid = 21'b000000001001111111011;
		14'b11001111111010:	sigmoid = 21'b000000001010000000101;
		14'b11001111111011:	sigmoid = 21'b000000001010000001111;
		14'b11001111111100:	sigmoid = 21'b000000001010000011001;
		14'b11001111111101:	sigmoid = 21'b000000001010000100011;
		14'b11001111111110:	sigmoid = 21'b000000001010000101101;
		14'b11001111111111:	sigmoid = 21'b000000001010000110111;
		14'b11010000000000:	sigmoid = 21'b000000001010001000001;
		14'b11010000000001:	sigmoid = 21'b000000001010001001011;
		14'b11010000000010:	sigmoid = 21'b000000001010001010101;
		14'b11010000000011:	sigmoid = 21'b000000001010001011111;
		14'b11010000000100:	sigmoid = 21'b000000001010001101010;
		14'b11010000000101:	sigmoid = 21'b000000001010001110100;
		14'b11010000000110:	sigmoid = 21'b000000001010001111110;
		14'b11010000000111:	sigmoid = 21'b000000001010010001000;
		14'b11010000001000:	sigmoid = 21'b000000001010010010010;
		14'b11010000001001:	sigmoid = 21'b000000001010010011101;
		14'b11010000001010:	sigmoid = 21'b000000001010010100111;
		14'b11010000001011:	sigmoid = 21'b000000001010010110001;
		14'b11010000001100:	sigmoid = 21'b000000001010010111100;
		14'b11010000001101:	sigmoid = 21'b000000001010011000110;
		14'b11010000001110:	sigmoid = 21'b000000001010011010000;
		14'b11010000001111:	sigmoid = 21'b000000001010011011011;
		14'b11010000010000:	sigmoid = 21'b000000001010011100101;
		14'b11010000010001:	sigmoid = 21'b000000001010011110000;
		14'b11010000010010:	sigmoid = 21'b000000001010011111010;
		14'b11010000010011:	sigmoid = 21'b000000001010100000101;
		14'b11010000010100:	sigmoid = 21'b000000001010100001111;
		14'b11010000010101:	sigmoid = 21'b000000001010100011010;
		14'b11010000010110:	sigmoid = 21'b000000001010100100100;
		14'b11010000010111:	sigmoid = 21'b000000001010100101111;
		14'b11010000011000:	sigmoid = 21'b000000001010100111001;
		14'b11010000011001:	sigmoid = 21'b000000001010101000100;
		14'b11010000011010:	sigmoid = 21'b000000001010101001110;
		14'b11010000011011:	sigmoid = 21'b000000001010101011001;
		14'b11010000011100:	sigmoid = 21'b000000001010101100100;
		14'b11010000011101:	sigmoid = 21'b000000001010101101110;
		14'b11010000011110:	sigmoid = 21'b000000001010101111001;
		14'b11010000011111:	sigmoid = 21'b000000001010110000100;
		14'b11010000100000:	sigmoid = 21'b000000001010110001111;
		14'b11010000100001:	sigmoid = 21'b000000001010110011001;
		14'b11010000100010:	sigmoid = 21'b000000001010110100100;
		14'b11010000100011:	sigmoid = 21'b000000001010110101111;
		14'b11010000100100:	sigmoid = 21'b000000001010110111010;
		14'b11010000100101:	sigmoid = 21'b000000001010111000101;
		14'b11010000100110:	sigmoid = 21'b000000001010111001111;
		14'b11010000100111:	sigmoid = 21'b000000001010111011010;
		14'b11010000101000:	sigmoid = 21'b000000001010111100101;
		14'b11010000101001:	sigmoid = 21'b000000001010111110000;
		14'b11010000101010:	sigmoid = 21'b000000001010111111011;
		14'b11010000101011:	sigmoid = 21'b000000001011000000110;
		14'b11010000101100:	sigmoid = 21'b000000001011000010001;
		14'b11010000101101:	sigmoid = 21'b000000001011000011100;
		14'b11010000101110:	sigmoid = 21'b000000001011000100111;
		14'b11010000101111:	sigmoid = 21'b000000001011000110010;
		14'b11010000110000:	sigmoid = 21'b000000001011000111101;
		14'b11010000110001:	sigmoid = 21'b000000001011001001000;
		14'b11010000110010:	sigmoid = 21'b000000001011001010011;
		14'b11010000110011:	sigmoid = 21'b000000001011001011111;
		14'b11010000110100:	sigmoid = 21'b000000001011001101010;
		14'b11010000110101:	sigmoid = 21'b000000001011001110101;
		14'b11010000110110:	sigmoid = 21'b000000001011010000000;
		14'b11010000110111:	sigmoid = 21'b000000001011010001011;
		14'b11010000111000:	sigmoid = 21'b000000001011010010111;
		14'b11010000111001:	sigmoid = 21'b000000001011010100010;
		14'b11010000111010:	sigmoid = 21'b000000001011010101101;
		14'b11010000111011:	sigmoid = 21'b000000001011010111001;
		14'b11010000111100:	sigmoid = 21'b000000001011011000100;
		14'b11010000111101:	sigmoid = 21'b000000001011011001111;
		14'b11010000111110:	sigmoid = 21'b000000001011011011011;
		14'b11010000111111:	sigmoid = 21'b000000001011011100110;
		14'b11010001000000:	sigmoid = 21'b000000001011011110001;
		14'b11010001000001:	sigmoid = 21'b000000001011011111101;
		14'b11010001000010:	sigmoid = 21'b000000001011100001000;
		14'b11010001000011:	sigmoid = 21'b000000001011100010100;
		14'b11010001000100:	sigmoid = 21'b000000001011100011111;
		14'b11010001000101:	sigmoid = 21'b000000001011100101011;
		14'b11010001000110:	sigmoid = 21'b000000001011100110111;
		14'b11010001000111:	sigmoid = 21'b000000001011101000010;
		14'b11010001001000:	sigmoid = 21'b000000001011101001110;
		14'b11010001001001:	sigmoid = 21'b000000001011101011001;
		14'b11010001001010:	sigmoid = 21'b000000001011101100101;
		14'b11010001001011:	sigmoid = 21'b000000001011101110001;
		14'b11010001001100:	sigmoid = 21'b000000001011101111100;
		14'b11010001001101:	sigmoid = 21'b000000001011110001000;
		14'b11010001001110:	sigmoid = 21'b000000001011110010100;
		14'b11010001001111:	sigmoid = 21'b000000001011110100000;
		14'b11010001010000:	sigmoid = 21'b000000001011110101011;
		14'b11010001010001:	sigmoid = 21'b000000001011110110111;
		14'b11010001010010:	sigmoid = 21'b000000001011111000011;
		14'b11010001010011:	sigmoid = 21'b000000001011111001111;
		14'b11010001010100:	sigmoid = 21'b000000001011111011011;
		14'b11010001010101:	sigmoid = 21'b000000001011111100111;
		14'b11010001010110:	sigmoid = 21'b000000001011111110011;
		14'b11010001010111:	sigmoid = 21'b000000001011111111111;
		14'b11010001011000:	sigmoid = 21'b000000001100000001011;
		14'b11010001011001:	sigmoid = 21'b000000001100000010111;
		14'b11010001011010:	sigmoid = 21'b000000001100000100011;
		14'b11010001011011:	sigmoid = 21'b000000001100000101111;
		14'b11010001011100:	sigmoid = 21'b000000001100000111011;
		14'b11010001011101:	sigmoid = 21'b000000001100001000111;
		14'b11010001011110:	sigmoid = 21'b000000001100001010011;
		14'b11010001011111:	sigmoid = 21'b000000001100001011111;
		14'b11010001100000:	sigmoid = 21'b000000001100001101011;
		14'b11010001100001:	sigmoid = 21'b000000001100001110111;
		14'b11010001100010:	sigmoid = 21'b000000001100010000100;
		14'b11010001100011:	sigmoid = 21'b000000001100010010000;
		14'b11010001100100:	sigmoid = 21'b000000001100010011100;
		14'b11010001100101:	sigmoid = 21'b000000001100010101000;
		14'b11010001100110:	sigmoid = 21'b000000001100010110101;
		14'b11010001100111:	sigmoid = 21'b000000001100011000001;
		14'b11010001101000:	sigmoid = 21'b000000001100011001101;
		14'b11010001101001:	sigmoid = 21'b000000001100011011010;
		14'b11010001101010:	sigmoid = 21'b000000001100011100110;
		14'b11010001101011:	sigmoid = 21'b000000001100011110011;
		14'b11010001101100:	sigmoid = 21'b000000001100011111111;
		14'b11010001101101:	sigmoid = 21'b000000001100100001011;
		14'b11010001101110:	sigmoid = 21'b000000001100100011000;
		14'b11010001101111:	sigmoid = 21'b000000001100100100100;
		14'b11010001110000:	sigmoid = 21'b000000001100100110001;
		14'b11010001110001:	sigmoid = 21'b000000001100100111110;
		14'b11010001110010:	sigmoid = 21'b000000001100101001010;
		14'b11010001110011:	sigmoid = 21'b000000001100101010111;
		14'b11010001110100:	sigmoid = 21'b000000001100101100011;
		14'b11010001110101:	sigmoid = 21'b000000001100101110000;
		14'b11010001110110:	sigmoid = 21'b000000001100101111101;
		14'b11010001110111:	sigmoid = 21'b000000001100110001010;
		14'b11010001111000:	sigmoid = 21'b000000001100110010110;
		14'b11010001111001:	sigmoid = 21'b000000001100110100011;
		14'b11010001111010:	sigmoid = 21'b000000001100110110000;
		14'b11010001111011:	sigmoid = 21'b000000001100110111101;
		14'b11010001111100:	sigmoid = 21'b000000001100111001001;
		14'b11010001111101:	sigmoid = 21'b000000001100111010110;
		14'b11010001111110:	sigmoid = 21'b000000001100111100011;
		14'b11010001111111:	sigmoid = 21'b000000001100111110000;
		14'b11010010000000:	sigmoid = 21'b000000001100111111101;
		14'b11010010000001:	sigmoid = 21'b000000001101000001010;
		14'b11010010000010:	sigmoid = 21'b000000001101000010111;
		14'b11010010000011:	sigmoid = 21'b000000001101000100100;
		14'b11010010000100:	sigmoid = 21'b000000001101000110001;
		14'b11010010000101:	sigmoid = 21'b000000001101000111110;
		14'b11010010000110:	sigmoid = 21'b000000001101001001011;
		14'b11010010000111:	sigmoid = 21'b000000001101001011000;
		14'b11010010001000:	sigmoid = 21'b000000001101001100110;
		14'b11010010001001:	sigmoid = 21'b000000001101001110011;
		14'b11010010001010:	sigmoid = 21'b000000001101010000000;
		14'b11010010001011:	sigmoid = 21'b000000001101010001101;
		14'b11010010001100:	sigmoid = 21'b000000001101010011010;
		14'b11010010001101:	sigmoid = 21'b000000001101010101000;
		14'b11010010001110:	sigmoid = 21'b000000001101010110101;
		14'b11010010001111:	sigmoid = 21'b000000001101011000010;
		14'b11010010010000:	sigmoid = 21'b000000001101011010000;
		14'b11010010010001:	sigmoid = 21'b000000001101011011101;
		14'b11010010010010:	sigmoid = 21'b000000001101011101010;
		14'b11010010010011:	sigmoid = 21'b000000001101011111000;
		14'b11010010010100:	sigmoid = 21'b000000001101100000101;
		14'b11010010010101:	sigmoid = 21'b000000001101100010011;
		14'b11010010010110:	sigmoid = 21'b000000001101100100000;
		14'b11010010010111:	sigmoid = 21'b000000001101100101110;
		14'b11010010011000:	sigmoid = 21'b000000001101100111011;
		14'b11010010011001:	sigmoid = 21'b000000001101101001001;
		14'b11010010011010:	sigmoid = 21'b000000001101101010111;
		14'b11010010011011:	sigmoid = 21'b000000001101101100100;
		14'b11010010011100:	sigmoid = 21'b000000001101101110010;
		14'b11010010011101:	sigmoid = 21'b000000001101110000000;
		14'b11010010011110:	sigmoid = 21'b000000001101110001101;
		14'b11010010011111:	sigmoid = 21'b000000001101110011011;
		14'b11010010100000:	sigmoid = 21'b000000001101110101001;
		14'b11010010100001:	sigmoid = 21'b000000001101110110111;
		14'b11010010100010:	sigmoid = 21'b000000001101111000100;
		14'b11010010100011:	sigmoid = 21'b000000001101111010010;
		14'b11010010100100:	sigmoid = 21'b000000001101111100000;
		14'b11010010100101:	sigmoid = 21'b000000001101111101110;
		14'b11010010100110:	sigmoid = 21'b000000001101111111100;
		14'b11010010100111:	sigmoid = 21'b000000001110000001010;
		14'b11010010101000:	sigmoid = 21'b000000001110000011000;
		14'b11010010101001:	sigmoid = 21'b000000001110000100110;
		14'b11010010101010:	sigmoid = 21'b000000001110000110100;
		14'b11010010101011:	sigmoid = 21'b000000001110001000010;
		14'b11010010101100:	sigmoid = 21'b000000001110001010000;
		14'b11010010101101:	sigmoid = 21'b000000001110001011110;
		14'b11010010101110:	sigmoid = 21'b000000001110001101100;
		14'b11010010101111:	sigmoid = 21'b000000001110001111011;
		14'b11010010110000:	sigmoid = 21'b000000001110010001001;
		14'b11010010110001:	sigmoid = 21'b000000001110010010111;
		14'b11010010110010:	sigmoid = 21'b000000001110010100101;
		14'b11010010110011:	sigmoid = 21'b000000001110010110100;
		14'b11010010110100:	sigmoid = 21'b000000001110011000010;
		14'b11010010110101:	sigmoid = 21'b000000001110011010000;
		14'b11010010110110:	sigmoid = 21'b000000001110011011111;
		14'b11010010110111:	sigmoid = 21'b000000001110011101101;
		14'b11010010111000:	sigmoid = 21'b000000001110011111011;
		14'b11010010111001:	sigmoid = 21'b000000001110100001010;
		14'b11010010111010:	sigmoid = 21'b000000001110100011000;
		14'b11010010111011:	sigmoid = 21'b000000001110100100111;
		14'b11010010111100:	sigmoid = 21'b000000001110100110101;
		14'b11010010111101:	sigmoid = 21'b000000001110101000100;
		14'b11010010111110:	sigmoid = 21'b000000001110101010011;
		14'b11010010111111:	sigmoid = 21'b000000001110101100001;
		14'b11010011000000:	sigmoid = 21'b000000001110101110000;
		14'b11010011000001:	sigmoid = 21'b000000001110101111111;
		14'b11010011000010:	sigmoid = 21'b000000001110110001101;
		14'b11010011000011:	sigmoid = 21'b000000001110110011100;
		14'b11010011000100:	sigmoid = 21'b000000001110110101011;
		14'b11010011000101:	sigmoid = 21'b000000001110110111010;
		14'b11010011000110:	sigmoid = 21'b000000001110111001000;
		14'b11010011000111:	sigmoid = 21'b000000001110111010111;
		14'b11010011001000:	sigmoid = 21'b000000001110111100110;
		14'b11010011001001:	sigmoid = 21'b000000001110111110101;
		14'b11010011001010:	sigmoid = 21'b000000001111000000100;
		14'b11010011001011:	sigmoid = 21'b000000001111000010011;
		14'b11010011001100:	sigmoid = 21'b000000001111000100010;
		14'b11010011001101:	sigmoid = 21'b000000001111000110001;
		14'b11010011001110:	sigmoid = 21'b000000001111001000000;
		14'b11010011001111:	sigmoid = 21'b000000001111001001111;
		14'b11010011010000:	sigmoid = 21'b000000001111001011110;
		14'b11010011010001:	sigmoid = 21'b000000001111001101101;
		14'b11010011010010:	sigmoid = 21'b000000001111001111100;
		14'b11010011010011:	sigmoid = 21'b000000001111010001100;
		14'b11010011010100:	sigmoid = 21'b000000001111010011011;
		14'b11010011010101:	sigmoid = 21'b000000001111010101010;
		14'b11010011010110:	sigmoid = 21'b000000001111010111001;
		14'b11010011010111:	sigmoid = 21'b000000001111011001001;
		14'b11010011011000:	sigmoid = 21'b000000001111011011000;
		14'b11010011011001:	sigmoid = 21'b000000001111011101000;
		14'b11010011011010:	sigmoid = 21'b000000001111011110111;
		14'b11010011011011:	sigmoid = 21'b000000001111100000110;
		14'b11010011011100:	sigmoid = 21'b000000001111100010110;
		14'b11010011011101:	sigmoid = 21'b000000001111100100101;
		14'b11010011011110:	sigmoid = 21'b000000001111100110101;
		14'b11010011011111:	sigmoid = 21'b000000001111101000100;
		14'b11010011100000:	sigmoid = 21'b000000001111101010100;
		14'b11010011100001:	sigmoid = 21'b000000001111101100100;
		14'b11010011100010:	sigmoid = 21'b000000001111101110011;
		14'b11010011100011:	sigmoid = 21'b000000001111110000011;
		14'b11010011100100:	sigmoid = 21'b000000001111110010011;
		14'b11010011100101:	sigmoid = 21'b000000001111110100010;
		14'b11010011100110:	sigmoid = 21'b000000001111110110010;
		14'b11010011100111:	sigmoid = 21'b000000001111111000010;
		14'b11010011101000:	sigmoid = 21'b000000001111111010010;
		14'b11010011101001:	sigmoid = 21'b000000001111111100010;
		14'b11010011101010:	sigmoid = 21'b000000001111111110010;
		14'b11010011101011:	sigmoid = 21'b000000010000000000010;
		14'b11010011101100:	sigmoid = 21'b000000010000000010001;
		14'b11010011101101:	sigmoid = 21'b000000010000000100001;
		14'b11010011101110:	sigmoid = 21'b000000010000000110001;
		14'b11010011101111:	sigmoid = 21'b000000010000001000010;
		14'b11010011110000:	sigmoid = 21'b000000010000001010010;
		14'b11010011110001:	sigmoid = 21'b000000010000001100010;
		14'b11010011110010:	sigmoid = 21'b000000010000001110010;
		14'b11010011110011:	sigmoid = 21'b000000010000010000010;
		14'b11010011110100:	sigmoid = 21'b000000010000010010010;
		14'b11010011110101:	sigmoid = 21'b000000010000010100010;
		14'b11010011110110:	sigmoid = 21'b000000010000010110011;
		14'b11010011110111:	sigmoid = 21'b000000010000011000011;
		14'b11010011111000:	sigmoid = 21'b000000010000011010011;
		14'b11010011111001:	sigmoid = 21'b000000010000011100100;
		14'b11010011111010:	sigmoid = 21'b000000010000011110100;
		14'b11010011111011:	sigmoid = 21'b000000010000100000101;
		14'b11010011111100:	sigmoid = 21'b000000010000100010101;
		14'b11010011111101:	sigmoid = 21'b000000010000100100110;
		14'b11010011111110:	sigmoid = 21'b000000010000100110110;
		14'b11010011111111:	sigmoid = 21'b000000010000101000111;
		14'b11010100000000:	sigmoid = 21'b000000010000101010111;
		14'b11010100000001:	sigmoid = 21'b000000010000101101000;
		14'b11010100000010:	sigmoid = 21'b000000010000101111000;
		14'b11010100000011:	sigmoid = 21'b000000010000110001001;
		14'b11010100000100:	sigmoid = 21'b000000010000110011010;
		14'b11010100000101:	sigmoid = 21'b000000010000110101011;
		14'b11010100000110:	sigmoid = 21'b000000010000110111011;
		14'b11010100000111:	sigmoid = 21'b000000010000111001100;
		14'b11010100001000:	sigmoid = 21'b000000010000111011101;
		14'b11010100001001:	sigmoid = 21'b000000010000111101110;
		14'b11010100001010:	sigmoid = 21'b000000010000111111111;
		14'b11010100001011:	sigmoid = 21'b000000010001000010000;
		14'b11010100001100:	sigmoid = 21'b000000010001000100001;
		14'b11010100001101:	sigmoid = 21'b000000010001000110010;
		14'b11010100001110:	sigmoid = 21'b000000010001001000011;
		14'b11010100001111:	sigmoid = 21'b000000010001001010100;
		14'b11010100010000:	sigmoid = 21'b000000010001001100101;
		14'b11010100010001:	sigmoid = 21'b000000010001001110110;
		14'b11010100010010:	sigmoid = 21'b000000010001010000111;
		14'b11010100010011:	sigmoid = 21'b000000010001010011001;
		14'b11010100010100:	sigmoid = 21'b000000010001010101010;
		14'b11010100010101:	sigmoid = 21'b000000010001010111011;
		14'b11010100010110:	sigmoid = 21'b000000010001011001100;
		14'b11010100010111:	sigmoid = 21'b000000010001011011110;
		14'b11010100011000:	sigmoid = 21'b000000010001011101111;
		14'b11010100011001:	sigmoid = 21'b000000010001100000000;
		14'b11010100011010:	sigmoid = 21'b000000010001100010010;
		14'b11010100011011:	sigmoid = 21'b000000010001100100011;
		14'b11010100011100:	sigmoid = 21'b000000010001100110101;
		14'b11010100011101:	sigmoid = 21'b000000010001101000110;
		14'b11010100011110:	sigmoid = 21'b000000010001101011000;
		14'b11010100011111:	sigmoid = 21'b000000010001101101010;
		14'b11010100100000:	sigmoid = 21'b000000010001101111011;
		14'b11010100100001:	sigmoid = 21'b000000010001110001101;
		14'b11010100100010:	sigmoid = 21'b000000010001110011111;
		14'b11010100100011:	sigmoid = 21'b000000010001110110000;
		14'b11010100100100:	sigmoid = 21'b000000010001111000010;
		14'b11010100100101:	sigmoid = 21'b000000010001111010100;
		14'b11010100100110:	sigmoid = 21'b000000010001111100110;
		14'b11010100100111:	sigmoid = 21'b000000010001111111000;
		14'b11010100101000:	sigmoid = 21'b000000010010000001010;
		14'b11010100101001:	sigmoid = 21'b000000010010000011100;
		14'b11010100101010:	sigmoid = 21'b000000010010000101110;
		14'b11010100101011:	sigmoid = 21'b000000010010001000000;
		14'b11010100101100:	sigmoid = 21'b000000010010001010010;
		14'b11010100101101:	sigmoid = 21'b000000010010001100100;
		14'b11010100101110:	sigmoid = 21'b000000010010001110110;
		14'b11010100101111:	sigmoid = 21'b000000010010010001000;
		14'b11010100110000:	sigmoid = 21'b000000010010010011010;
		14'b11010100110001:	sigmoid = 21'b000000010010010101101;
		14'b11010100110010:	sigmoid = 21'b000000010010010111111;
		14'b11010100110011:	sigmoid = 21'b000000010010011010001;
		14'b11010100110100:	sigmoid = 21'b000000010010011100100;
		14'b11010100110101:	sigmoid = 21'b000000010010011110110;
		14'b11010100110110:	sigmoid = 21'b000000010010100001000;
		14'b11010100110111:	sigmoid = 21'b000000010010100011011;
		14'b11010100111000:	sigmoid = 21'b000000010010100101101;
		14'b11010100111001:	sigmoid = 21'b000000010010101000000;
		14'b11010100111010:	sigmoid = 21'b000000010010101010010;
		14'b11010100111011:	sigmoid = 21'b000000010010101100101;
		14'b11010100111100:	sigmoid = 21'b000000010010101111000;
		14'b11010100111101:	sigmoid = 21'b000000010010110001010;
		14'b11010100111110:	sigmoid = 21'b000000010010110011101;
		14'b11010100111111:	sigmoid = 21'b000000010010110110000;
		14'b11010101000000:	sigmoid = 21'b000000010010111000010;
		14'b11010101000001:	sigmoid = 21'b000000010010111010101;
		14'b11010101000010:	sigmoid = 21'b000000010010111101000;
		14'b11010101000011:	sigmoid = 21'b000000010010111111011;
		14'b11010101000100:	sigmoid = 21'b000000010011000001110;
		14'b11010101000101:	sigmoid = 21'b000000010011000100001;
		14'b11010101000110:	sigmoid = 21'b000000010011000110100;
		14'b11010101000111:	sigmoid = 21'b000000010011001000111;
		14'b11010101001000:	sigmoid = 21'b000000010011001011010;
		14'b11010101001001:	sigmoid = 21'b000000010011001101101;
		14'b11010101001010:	sigmoid = 21'b000000010011010000000;
		14'b11010101001011:	sigmoid = 21'b000000010011010010011;
		14'b11010101001100:	sigmoid = 21'b000000010011010100111;
		14'b11010101001101:	sigmoid = 21'b000000010011010111010;
		14'b11010101001110:	sigmoid = 21'b000000010011011001101;
		14'b11010101001111:	sigmoid = 21'b000000010011011100001;
		14'b11010101010000:	sigmoid = 21'b000000010011011110100;
		14'b11010101010001:	sigmoid = 21'b000000010011100000111;
		14'b11010101010010:	sigmoid = 21'b000000010011100011011;
		14'b11010101010011:	sigmoid = 21'b000000010011100101110;
		14'b11010101010100:	sigmoid = 21'b000000010011101000010;
		14'b11010101010101:	sigmoid = 21'b000000010011101010101;
		14'b11010101010110:	sigmoid = 21'b000000010011101101001;
		14'b11010101010111:	sigmoid = 21'b000000010011101111100;
		14'b11010101011000:	sigmoid = 21'b000000010011110010000;
		14'b11010101011001:	sigmoid = 21'b000000010011110100100;
		14'b11010101011010:	sigmoid = 21'b000000010011110111000;
		14'b11010101011011:	sigmoid = 21'b000000010011111001011;
		14'b11010101011100:	sigmoid = 21'b000000010011111011111;
		14'b11010101011101:	sigmoid = 21'b000000010011111110011;
		14'b11010101011110:	sigmoid = 21'b000000010100000000111;
		14'b11010101011111:	sigmoid = 21'b000000010100000011011;
		14'b11010101100000:	sigmoid = 21'b000000010100000101111;
		14'b11010101100001:	sigmoid = 21'b000000010100001000011;
		14'b11010101100010:	sigmoid = 21'b000000010100001010111;
		14'b11010101100011:	sigmoid = 21'b000000010100001101011;
		14'b11010101100100:	sigmoid = 21'b000000010100001111111;
		14'b11010101100101:	sigmoid = 21'b000000010100010010011;
		14'b11010101100110:	sigmoid = 21'b000000010100010101000;
		14'b11010101100111:	sigmoid = 21'b000000010100010111100;
		14'b11010101101000:	sigmoid = 21'b000000010100011010000;
		14'b11010101101001:	sigmoid = 21'b000000010100011100100;
		14'b11010101101010:	sigmoid = 21'b000000010100011111001;
		14'b11010101101011:	sigmoid = 21'b000000010100100001101;
		14'b11010101101100:	sigmoid = 21'b000000010100100100010;
		14'b11010101101101:	sigmoid = 21'b000000010100100110110;
		14'b11010101101110:	sigmoid = 21'b000000010100101001011;
		14'b11010101101111:	sigmoid = 21'b000000010100101011111;
		14'b11010101110000:	sigmoid = 21'b000000010100101110100;
		14'b11010101110001:	sigmoid = 21'b000000010100110001000;
		14'b11010101110010:	sigmoid = 21'b000000010100110011101;
		14'b11010101110011:	sigmoid = 21'b000000010100110110010;
		14'b11010101110100:	sigmoid = 21'b000000010100111000111;
		14'b11010101110101:	sigmoid = 21'b000000010100111011011;
		14'b11010101110110:	sigmoid = 21'b000000010100111110000;
		14'b11010101110111:	sigmoid = 21'b000000010101000000101;
		14'b11010101111000:	sigmoid = 21'b000000010101000011010;
		14'b11010101111001:	sigmoid = 21'b000000010101000101111;
		14'b11010101111010:	sigmoid = 21'b000000010101001000100;
		14'b11010101111011:	sigmoid = 21'b000000010101001011001;
		14'b11010101111100:	sigmoid = 21'b000000010101001101110;
		14'b11010101111101:	sigmoid = 21'b000000010101010000011;
		14'b11010101111110:	sigmoid = 21'b000000010101010011000;
		14'b11010101111111:	sigmoid = 21'b000000010101010101110;
		14'b11010110000000:	sigmoid = 21'b000000010101011000011;
		14'b11010110000001:	sigmoid = 21'b000000010101011011000;
		14'b11010110000010:	sigmoid = 21'b000000010101011101110;
		14'b11010110000011:	sigmoid = 21'b000000010101100000011;
		14'b11010110000100:	sigmoid = 21'b000000010101100011000;
		14'b11010110000101:	sigmoid = 21'b000000010101100101110;
		14'b11010110000110:	sigmoid = 21'b000000010101101000011;
		14'b11010110000111:	sigmoid = 21'b000000010101101011001;
		14'b11010110001000:	sigmoid = 21'b000000010101101101110;
		14'b11010110001001:	sigmoid = 21'b000000010101110000100;
		14'b11010110001010:	sigmoid = 21'b000000010101110011010;
		14'b11010110001011:	sigmoid = 21'b000000010101110101111;
		14'b11010110001100:	sigmoid = 21'b000000010101111000101;
		14'b11010110001101:	sigmoid = 21'b000000010101111011011;
		14'b11010110001110:	sigmoid = 21'b000000010101111110001;
		14'b11010110001111:	sigmoid = 21'b000000010110000000111;
		14'b11010110010000:	sigmoid = 21'b000000010110000011101;
		14'b11010110010001:	sigmoid = 21'b000000010110000110010;
		14'b11010110010010:	sigmoid = 21'b000000010110001001000;
		14'b11010110010011:	sigmoid = 21'b000000010110001011111;
		14'b11010110010100:	sigmoid = 21'b000000010110001110101;
		14'b11010110010101:	sigmoid = 21'b000000010110010001011;
		14'b11010110010110:	sigmoid = 21'b000000010110010100001;
		14'b11010110010111:	sigmoid = 21'b000000010110010110111;
		14'b11010110011000:	sigmoid = 21'b000000010110011001101;
		14'b11010110011001:	sigmoid = 21'b000000010110011100100;
		14'b11010110011010:	sigmoid = 21'b000000010110011111010;
		14'b11010110011011:	sigmoid = 21'b000000010110100010000;
		14'b11010110011100:	sigmoid = 21'b000000010110100100111;
		14'b11010110011101:	sigmoid = 21'b000000010110100111101;
		14'b11010110011110:	sigmoid = 21'b000000010110101010100;
		14'b11010110011111:	sigmoid = 21'b000000010110101101010;
		14'b11010110100000:	sigmoid = 21'b000000010110110000001;
		14'b11010110100001:	sigmoid = 21'b000000010110110011000;
		14'b11010110100010:	sigmoid = 21'b000000010110110101110;
		14'b11010110100011:	sigmoid = 21'b000000010110111000101;
		14'b11010110100100:	sigmoid = 21'b000000010110111011100;
		14'b11010110100101:	sigmoid = 21'b000000010110111110011;
		14'b11010110100110:	sigmoid = 21'b000000010111000001010;
		14'b11010110100111:	sigmoid = 21'b000000010111000100000;
		14'b11010110101000:	sigmoid = 21'b000000010111000110111;
		14'b11010110101001:	sigmoid = 21'b000000010111001001110;
		14'b11010110101010:	sigmoid = 21'b000000010111001100101;
		14'b11010110101011:	sigmoid = 21'b000000010111001111101;
		14'b11010110101100:	sigmoid = 21'b000000010111010010100;
		14'b11010110101101:	sigmoid = 21'b000000010111010101011;
		14'b11010110101110:	sigmoid = 21'b000000010111011000010;
		14'b11010110101111:	sigmoid = 21'b000000010111011011001;
		14'b11010110110000:	sigmoid = 21'b000000010111011110001;
		14'b11010110110001:	sigmoid = 21'b000000010111100001000;
		14'b11010110110010:	sigmoid = 21'b000000010111100011111;
		14'b11010110110011:	sigmoid = 21'b000000010111100110111;
		14'b11010110110100:	sigmoid = 21'b000000010111101001110;
		14'b11010110110101:	sigmoid = 21'b000000010111101100110;
		14'b11010110110110:	sigmoid = 21'b000000010111101111110;
		14'b11010110110111:	sigmoid = 21'b000000010111110010101;
		14'b11010110111000:	sigmoid = 21'b000000010111110101101;
		14'b11010110111001:	sigmoid = 21'b000000010111111000101;
		14'b11010110111010:	sigmoid = 21'b000000010111111011100;
		14'b11010110111011:	sigmoid = 21'b000000010111111110100;
		14'b11010110111100:	sigmoid = 21'b000000011000000001100;
		14'b11010110111101:	sigmoid = 21'b000000011000000100100;
		14'b11010110111110:	sigmoid = 21'b000000011000000111100;
		14'b11010110111111:	sigmoid = 21'b000000011000001010100;
		14'b11010111000000:	sigmoid = 21'b000000011000001101100;
		14'b11010111000001:	sigmoid = 21'b000000011000010000100;
		14'b11010111000010:	sigmoid = 21'b000000011000010011100;
		14'b11010111000011:	sigmoid = 21'b000000011000010110100;
		14'b11010111000100:	sigmoid = 21'b000000011000011001101;
		14'b11010111000101:	sigmoid = 21'b000000011000011100101;
		14'b11010111000110:	sigmoid = 21'b000000011000011111101;
		14'b11010111000111:	sigmoid = 21'b000000011000100010110;
		14'b11010111001000:	sigmoid = 21'b000000011000100101110;
		14'b11010111001001:	sigmoid = 21'b000000011000101000110;
		14'b11010111001010:	sigmoid = 21'b000000011000101011111;
		14'b11010111001011:	sigmoid = 21'b000000011000101110111;
		14'b11010111001100:	sigmoid = 21'b000000011000110010000;
		14'b11010111001101:	sigmoid = 21'b000000011000110101001;
		14'b11010111001110:	sigmoid = 21'b000000011000111000001;
		14'b11010111001111:	sigmoid = 21'b000000011000111011010;
		14'b11010111010000:	sigmoid = 21'b000000011000111110011;
		14'b11010111010001:	sigmoid = 21'b000000011001000001100;
		14'b11010111010010:	sigmoid = 21'b000000011001000100101;
		14'b11010111010011:	sigmoid = 21'b000000011001000111110;
		14'b11010111010100:	sigmoid = 21'b000000011001001010111;
		14'b11010111010101:	sigmoid = 21'b000000011001001110000;
		14'b11010111010110:	sigmoid = 21'b000000011001010001001;
		14'b11010111010111:	sigmoid = 21'b000000011001010100010;
		14'b11010111011000:	sigmoid = 21'b000000011001010111011;
		14'b11010111011001:	sigmoid = 21'b000000011001011010100;
		14'b11010111011010:	sigmoid = 21'b000000011001011101110;
		14'b11010111011011:	sigmoid = 21'b000000011001100000111;
		14'b11010111011100:	sigmoid = 21'b000000011001100100000;
		14'b11010111011101:	sigmoid = 21'b000000011001100111010;
		14'b11010111011110:	sigmoid = 21'b000000011001101010011;
		14'b11010111011111:	sigmoid = 21'b000000011001101101101;
		14'b11010111100000:	sigmoid = 21'b000000011001110000110;
		14'b11010111100001:	sigmoid = 21'b000000011001110100000;
		14'b11010111100010:	sigmoid = 21'b000000011001110111010;
		14'b11010111100011:	sigmoid = 21'b000000011001111010011;
		14'b11010111100100:	sigmoid = 21'b000000011001111101101;
		14'b11010111100101:	sigmoid = 21'b000000011010000000111;
		14'b11010111100110:	sigmoid = 21'b000000011010000100001;
		14'b11010111100111:	sigmoid = 21'b000000011010000111011;
		14'b11010111101000:	sigmoid = 21'b000000011010001010101;
		14'b11010111101001:	sigmoid = 21'b000000011010001101111;
		14'b11010111101010:	sigmoid = 21'b000000011010010001001;
		14'b11010111101011:	sigmoid = 21'b000000011010010100011;
		14'b11010111101100:	sigmoid = 21'b000000011010010111101;
		14'b11010111101101:	sigmoid = 21'b000000011010011010111;
		14'b11010111101110:	sigmoid = 21'b000000011010011110010;
		14'b11010111101111:	sigmoid = 21'b000000011010100001100;
		14'b11010111110000:	sigmoid = 21'b000000011010100100110;
		14'b11010111110001:	sigmoid = 21'b000000011010101000001;
		14'b11010111110010:	sigmoid = 21'b000000011010101011011;
		14'b11010111110011:	sigmoid = 21'b000000011010101110110;
		14'b11010111110100:	sigmoid = 21'b000000011010110010000;
		14'b11010111110101:	sigmoid = 21'b000000011010110101011;
		14'b11010111110110:	sigmoid = 21'b000000011010111000110;
		14'b11010111110111:	sigmoid = 21'b000000011010111100000;
		14'b11010111111000:	sigmoid = 21'b000000011010111111011;
		14'b11010111111001:	sigmoid = 21'b000000011011000010110;
		14'b11010111111010:	sigmoid = 21'b000000011011000110001;
		14'b11010111111011:	sigmoid = 21'b000000011011001001100;
		14'b11010111111100:	sigmoid = 21'b000000011011001100111;
		14'b11010111111101:	sigmoid = 21'b000000011011010000010;
		14'b11010111111110:	sigmoid = 21'b000000011011010011101;
		14'b11010111111111:	sigmoid = 21'b000000011011010111000;
		14'b11011000000000:	sigmoid = 21'b000000011011011010011;
		14'b11011000000001:	sigmoid = 21'b000000011011011101111;
		14'b11011000000010:	sigmoid = 21'b000000011011100001010;
		14'b11011000000011:	sigmoid = 21'b000000011011100100101;
		14'b11011000000100:	sigmoid = 21'b000000011011101000001;
		14'b11011000000101:	sigmoid = 21'b000000011011101011100;
		14'b11011000000110:	sigmoid = 21'b000000011011101111000;
		14'b11011000000111:	sigmoid = 21'b000000011011110010011;
		14'b11011000001000:	sigmoid = 21'b000000011011110101111;
		14'b11011000001001:	sigmoid = 21'b000000011011111001011;
		14'b11011000001010:	sigmoid = 21'b000000011011111100110;
		14'b11011000001011:	sigmoid = 21'b000000011100000000010;
		14'b11011000001100:	sigmoid = 21'b000000011100000011110;
		14'b11011000001101:	sigmoid = 21'b000000011100000111010;
		14'b11011000001110:	sigmoid = 21'b000000011100001010110;
		14'b11011000001111:	sigmoid = 21'b000000011100001110010;
		14'b11011000010000:	sigmoid = 21'b000000011100010001110;
		14'b11011000010001:	sigmoid = 21'b000000011100010101010;
		14'b11011000010010:	sigmoid = 21'b000000011100011000110;
		14'b11011000010011:	sigmoid = 21'b000000011100011100010;
		14'b11011000010100:	sigmoid = 21'b000000011100011111111;
		14'b11011000010101:	sigmoid = 21'b000000011100100011011;
		14'b11011000010110:	sigmoid = 21'b000000011100100110111;
		14'b11011000010111:	sigmoid = 21'b000000011100101010100;
		14'b11011000011000:	sigmoid = 21'b000000011100101110000;
		14'b11011000011001:	sigmoid = 21'b000000011100110001101;
		14'b11011000011010:	sigmoid = 21'b000000011100110101001;
		14'b11011000011011:	sigmoid = 21'b000000011100111000110;
		14'b11011000011100:	sigmoid = 21'b000000011100111100011;
		14'b11011000011101:	sigmoid = 21'b000000011101000000000;
		14'b11011000011110:	sigmoid = 21'b000000011101000011100;
		14'b11011000011111:	sigmoid = 21'b000000011101000111001;
		14'b11011000100000:	sigmoid = 21'b000000011101001010110;
		14'b11011000100001:	sigmoid = 21'b000000011101001110011;
		14'b11011000100010:	sigmoid = 21'b000000011101010010000;
		14'b11011000100011:	sigmoid = 21'b000000011101010101101;
		14'b11011000100100:	sigmoid = 21'b000000011101011001011;
		14'b11011000100101:	sigmoid = 21'b000000011101011101000;
		14'b11011000100110:	sigmoid = 21'b000000011101100000101;
		14'b11011000100111:	sigmoid = 21'b000000011101100100010;
		14'b11011000101000:	sigmoid = 21'b000000011101101000000;
		14'b11011000101001:	sigmoid = 21'b000000011101101011101;
		14'b11011000101010:	sigmoid = 21'b000000011101101111011;
		14'b11011000101011:	sigmoid = 21'b000000011101110011000;
		14'b11011000101100:	sigmoid = 21'b000000011101110110110;
		14'b11011000101101:	sigmoid = 21'b000000011101111010011;
		14'b11011000101110:	sigmoid = 21'b000000011101111110001;
		14'b11011000101111:	sigmoid = 21'b000000011110000001111;
		14'b11011000110000:	sigmoid = 21'b000000011110000101101;
		14'b11011000110001:	sigmoid = 21'b000000011110001001011;
		14'b11011000110010:	sigmoid = 21'b000000011110001101001;
		14'b11011000110011:	sigmoid = 21'b000000011110010000111;
		14'b11011000110100:	sigmoid = 21'b000000011110010100101;
		14'b11011000110101:	sigmoid = 21'b000000011110011000011;
		14'b11011000110110:	sigmoid = 21'b000000011110011100001;
		14'b11011000110111:	sigmoid = 21'b000000011110011111111;
		14'b11011000111000:	sigmoid = 21'b000000011110100011110;
		14'b11011000111001:	sigmoid = 21'b000000011110100111100;
		14'b11011000111010:	sigmoid = 21'b000000011110101011010;
		14'b11011000111011:	sigmoid = 21'b000000011110101111001;
		14'b11011000111100:	sigmoid = 21'b000000011110110010111;
		14'b11011000111101:	sigmoid = 21'b000000011110110110110;
		14'b11011000111110:	sigmoid = 21'b000000011110111010101;
		14'b11011000111111:	sigmoid = 21'b000000011110111110011;
		14'b11011001000000:	sigmoid = 21'b000000011111000010010;
		14'b11011001000001:	sigmoid = 21'b000000011111000110001;
		14'b11011001000010:	sigmoid = 21'b000000011111001010000;
		14'b11011001000011:	sigmoid = 21'b000000011111001101111;
		14'b11011001000100:	sigmoid = 21'b000000011111010001110;
		14'b11011001000101:	sigmoid = 21'b000000011111010101101;
		14'b11011001000110:	sigmoid = 21'b000000011111011001100;
		14'b11011001000111:	sigmoid = 21'b000000011111011101011;
		14'b11011001001000:	sigmoid = 21'b000000011111100001010;
		14'b11011001001001:	sigmoid = 21'b000000011111100101010;
		14'b11011001001010:	sigmoid = 21'b000000011111101001001;
		14'b11011001001011:	sigmoid = 21'b000000011111101101001;
		14'b11011001001100:	sigmoid = 21'b000000011111110001000;
		14'b11011001001101:	sigmoid = 21'b000000011111110101000;
		14'b11011001001110:	sigmoid = 21'b000000011111111000111;
		14'b11011001001111:	sigmoid = 21'b000000011111111100111;
		14'b11011001010000:	sigmoid = 21'b000000100000000000111;
		14'b11011001010001:	sigmoid = 21'b000000100000000100110;
		14'b11011001010010:	sigmoid = 21'b000000100000001000110;
		14'b11011001010011:	sigmoid = 21'b000000100000001100110;
		14'b11011001010100:	sigmoid = 21'b000000100000010000110;
		14'b11011001010101:	sigmoid = 21'b000000100000010100110;
		14'b11011001010110:	sigmoid = 21'b000000100000011000110;
		14'b11011001010111:	sigmoid = 21'b000000100000011100110;
		14'b11011001011000:	sigmoid = 21'b000000100000100000111;
		14'b11011001011001:	sigmoid = 21'b000000100000100100111;
		14'b11011001011010:	sigmoid = 21'b000000100000101000111;
		14'b11011001011011:	sigmoid = 21'b000000100000101101000;
		14'b11011001011100:	sigmoid = 21'b000000100000110001000;
		14'b11011001011101:	sigmoid = 21'b000000100000110101001;
		14'b11011001011110:	sigmoid = 21'b000000100000111001001;
		14'b11011001011111:	sigmoid = 21'b000000100000111101010;
		14'b11011001100000:	sigmoid = 21'b000000100001000001011;
		14'b11011001100001:	sigmoid = 21'b000000100001000101100;
		14'b11011001100010:	sigmoid = 21'b000000100001001001100;
		14'b11011001100011:	sigmoid = 21'b000000100001001101101;
		14'b11011001100100:	sigmoid = 21'b000000100001010001110;
		14'b11011001100101:	sigmoid = 21'b000000100001010101111;
		14'b11011001100110:	sigmoid = 21'b000000100001011010000;
		14'b11011001100111:	sigmoid = 21'b000000100001011110010;
		14'b11011001101000:	sigmoid = 21'b000000100001100010011;
		14'b11011001101001:	sigmoid = 21'b000000100001100110100;
		14'b11011001101010:	sigmoid = 21'b000000100001101010101;
		14'b11011001101011:	sigmoid = 21'b000000100001101110111;
		14'b11011001101100:	sigmoid = 21'b000000100001110011000;
		14'b11011001101101:	sigmoid = 21'b000000100001110111010;
		14'b11011001101110:	sigmoid = 21'b000000100001111011100;
		14'b11011001101111:	sigmoid = 21'b000000100001111111101;
		14'b11011001110000:	sigmoid = 21'b000000100010000011111;
		14'b11011001110001:	sigmoid = 21'b000000100010001000001;
		14'b11011001110010:	sigmoid = 21'b000000100010001100011;
		14'b11011001110011:	sigmoid = 21'b000000100010010000101;
		14'b11011001110100:	sigmoid = 21'b000000100010010100111;
		14'b11011001110101:	sigmoid = 21'b000000100010011001001;
		14'b11011001110110:	sigmoid = 21'b000000100010011101011;
		14'b11011001110111:	sigmoid = 21'b000000100010100001101;
		14'b11011001111000:	sigmoid = 21'b000000100010100101111;
		14'b11011001111001:	sigmoid = 21'b000000100010101010010;
		14'b11011001111010:	sigmoid = 21'b000000100010101110100;
		14'b11011001111011:	sigmoid = 21'b000000100010110010110;
		14'b11011001111100:	sigmoid = 21'b000000100010110111001;
		14'b11011001111101:	sigmoid = 21'b000000100010111011100;
		14'b11011001111110:	sigmoid = 21'b000000100010111111110;
		14'b11011001111111:	sigmoid = 21'b000000100011000100001;
		14'b11011010000000:	sigmoid = 21'b000000100011001000100;
		14'b11011010000001:	sigmoid = 21'b000000100011001100111;
		14'b11011010000010:	sigmoid = 21'b000000100011010001010;
		14'b11011010000011:	sigmoid = 21'b000000100011010101101;
		14'b11011010000100:	sigmoid = 21'b000000100011011010000;
		14'b11011010000101:	sigmoid = 21'b000000100011011110011;
		14'b11011010000110:	sigmoid = 21'b000000100011100010110;
		14'b11011010000111:	sigmoid = 21'b000000100011100111001;
		14'b11011010001000:	sigmoid = 21'b000000100011101011101;
		14'b11011010001001:	sigmoid = 21'b000000100011110000000;
		14'b11011010001010:	sigmoid = 21'b000000100011110100011;
		14'b11011010001011:	sigmoid = 21'b000000100011111000111;
		14'b11011010001100:	sigmoid = 21'b000000100011111101011;
		14'b11011010001101:	sigmoid = 21'b000000100100000001110;
		14'b11011010001110:	sigmoid = 21'b000000100100000110010;
		14'b11011010001111:	sigmoid = 21'b000000100100001010110;
		14'b11011010010000:	sigmoid = 21'b000000100100001111010;
		14'b11011010010001:	sigmoid = 21'b000000100100010011110;
		14'b11011010010010:	sigmoid = 21'b000000100100011000010;
		14'b11011010010011:	sigmoid = 21'b000000100100011100110;
		14'b11011010010100:	sigmoid = 21'b000000100100100001010;
		14'b11011010010101:	sigmoid = 21'b000000100100100101110;
		14'b11011010010110:	sigmoid = 21'b000000100100101010011;
		14'b11011010010111:	sigmoid = 21'b000000100100101110111;
		14'b11011010011000:	sigmoid = 21'b000000100100110011011;
		14'b11011010011001:	sigmoid = 21'b000000100100111000000;
		14'b11011010011010:	sigmoid = 21'b000000100100111100100;
		14'b11011010011011:	sigmoid = 21'b000000100101000001001;
		14'b11011010011100:	sigmoid = 21'b000000100101000101110;
		14'b11011010011101:	sigmoid = 21'b000000100101001010011;
		14'b11011010011110:	sigmoid = 21'b000000100101001110111;
		14'b11011010011111:	sigmoid = 21'b000000100101010011100;
		14'b11011010100000:	sigmoid = 21'b000000100101011000001;
		14'b11011010100001:	sigmoid = 21'b000000100101011100110;
		14'b11011010100010:	sigmoid = 21'b000000100101100001100;
		14'b11011010100011:	sigmoid = 21'b000000100101100110001;
		14'b11011010100100:	sigmoid = 21'b000000100101101010110;
		14'b11011010100101:	sigmoid = 21'b000000100101101111011;
		14'b11011010100110:	sigmoid = 21'b000000100101110100001;
		14'b11011010100111:	sigmoid = 21'b000000100101111000110;
		14'b11011010101000:	sigmoid = 21'b000000100101111101100;
		14'b11011010101001:	sigmoid = 21'b000000100110000010010;
		14'b11011010101010:	sigmoid = 21'b000000100110000110111;
		14'b11011010101011:	sigmoid = 21'b000000100110001011101;
		14'b11011010101100:	sigmoid = 21'b000000100110010000011;
		14'b11011010101101:	sigmoid = 21'b000000100110010101001;
		14'b11011010101110:	sigmoid = 21'b000000100110011001111;
		14'b11011010101111:	sigmoid = 21'b000000100110011110101;
		14'b11011010110000:	sigmoid = 21'b000000100110100011011;
		14'b11011010110001:	sigmoid = 21'b000000100110101000001;
		14'b11011010110010:	sigmoid = 21'b000000100110101101000;
		14'b11011010110011:	sigmoid = 21'b000000100110110001110;
		14'b11011010110100:	sigmoid = 21'b000000100110110110100;
		14'b11011010110101:	sigmoid = 21'b000000100110111011011;
		14'b11011010110110:	sigmoid = 21'b000000100111000000010;
		14'b11011010110111:	sigmoid = 21'b000000100111000101000;
		14'b11011010111000:	sigmoid = 21'b000000100111001001111;
		14'b11011010111001:	sigmoid = 21'b000000100111001110110;
		14'b11011010111010:	sigmoid = 21'b000000100111010011101;
		14'b11011010111011:	sigmoid = 21'b000000100111011000100;
		14'b11011010111100:	sigmoid = 21'b000000100111011101011;
		14'b11011010111101:	sigmoid = 21'b000000100111100010010;
		14'b11011010111110:	sigmoid = 21'b000000100111100111001;
		14'b11011010111111:	sigmoid = 21'b000000100111101100000;
		14'b11011011000000:	sigmoid = 21'b000000100111110001000;
		14'b11011011000001:	sigmoid = 21'b000000100111110101111;
		14'b11011011000010:	sigmoid = 21'b000000100111111010111;
		14'b11011011000011:	sigmoid = 21'b000000100111111111110;
		14'b11011011000100:	sigmoid = 21'b000000101000000100110;
		14'b11011011000101:	sigmoid = 21'b000000101000001001101;
		14'b11011011000110:	sigmoid = 21'b000000101000001110101;
		14'b11011011000111:	sigmoid = 21'b000000101000010011101;
		14'b11011011001000:	sigmoid = 21'b000000101000011000101;
		14'b11011011001001:	sigmoid = 21'b000000101000011101101;
		14'b11011011001010:	sigmoid = 21'b000000101000100010101;
		14'b11011011001011:	sigmoid = 21'b000000101000100111101;
		14'b11011011001100:	sigmoid = 21'b000000101000101100110;
		14'b11011011001101:	sigmoid = 21'b000000101000110001110;
		14'b11011011001110:	sigmoid = 21'b000000101000110110110;
		14'b11011011001111:	sigmoid = 21'b000000101000111011111;
		14'b11011011010000:	sigmoid = 21'b000000101001000000111;
		14'b11011011010001:	sigmoid = 21'b000000101001000110000;
		14'b11011011010010:	sigmoid = 21'b000000101001001011001;
		14'b11011011010011:	sigmoid = 21'b000000101001010000010;
		14'b11011011010100:	sigmoid = 21'b000000101001010101011;
		14'b11011011010101:	sigmoid = 21'b000000101001011010011;
		14'b11011011010110:	sigmoid = 21'b000000101001011111101;
		14'b11011011010111:	sigmoid = 21'b000000101001100100110;
		14'b11011011011000:	sigmoid = 21'b000000101001101001111;
		14'b11011011011001:	sigmoid = 21'b000000101001101111000;
		14'b11011011011010:	sigmoid = 21'b000000101001110100001;
		14'b11011011011011:	sigmoid = 21'b000000101001111001011;
		14'b11011011011100:	sigmoid = 21'b000000101001111110100;
		14'b11011011011101:	sigmoid = 21'b000000101010000011110;
		14'b11011011011110:	sigmoid = 21'b000000101010001001000;
		14'b11011011011111:	sigmoid = 21'b000000101010001110001;
		14'b11011011100000:	sigmoid = 21'b000000101010010011011;
		14'b11011011100001:	sigmoid = 21'b000000101010011000101;
		14'b11011011100010:	sigmoid = 21'b000000101010011101111;
		14'b11011011100011:	sigmoid = 21'b000000101010100011001;
		14'b11011011100100:	sigmoid = 21'b000000101010101000011;
		14'b11011011100101:	sigmoid = 21'b000000101010101101110;
		14'b11011011100110:	sigmoid = 21'b000000101010110011000;
		14'b11011011100111:	sigmoid = 21'b000000101010111000010;
		14'b11011011101000:	sigmoid = 21'b000000101010111101101;
		14'b11011011101001:	sigmoid = 21'b000000101011000010111;
		14'b11011011101010:	sigmoid = 21'b000000101011001000010;
		14'b11011011101011:	sigmoid = 21'b000000101011001101101;
		14'b11011011101100:	sigmoid = 21'b000000101011010010111;
		14'b11011011101101:	sigmoid = 21'b000000101011011000010;
		14'b11011011101110:	sigmoid = 21'b000000101011011101101;
		14'b11011011101111:	sigmoid = 21'b000000101011100011000;
		14'b11011011110000:	sigmoid = 21'b000000101011101000011;
		14'b11011011110001:	sigmoid = 21'b000000101011101101111;
		14'b11011011110010:	sigmoid = 21'b000000101011110011010;
		14'b11011011110011:	sigmoid = 21'b000000101011111000101;
		14'b11011011110100:	sigmoid = 21'b000000101011111110001;
		14'b11011011110101:	sigmoid = 21'b000000101100000011100;
		14'b11011011110110:	sigmoid = 21'b000000101100001001000;
		14'b11011011110111:	sigmoid = 21'b000000101100001110100;
		14'b11011011111000:	sigmoid = 21'b000000101100010011111;
		14'b11011011111001:	sigmoid = 21'b000000101100011001011;
		14'b11011011111010:	sigmoid = 21'b000000101100011110111;
		14'b11011011111011:	sigmoid = 21'b000000101100100100011;
		14'b11011011111100:	sigmoid = 21'b000000101100101001111;
		14'b11011011111101:	sigmoid = 21'b000000101100101111100;
		14'b11011011111110:	sigmoid = 21'b000000101100110101000;
		14'b11011011111111:	sigmoid = 21'b000000101100111010100;
		14'b11011100000000:	sigmoid = 21'b000000101101000000001;
		14'b11011100000001:	sigmoid = 21'b000000101101000101101;
		14'b11011100000010:	sigmoid = 21'b000000101101001011010;
		14'b11011100000011:	sigmoid = 21'b000000101101010000111;
		14'b11011100000100:	sigmoid = 21'b000000101101010110100;
		14'b11011100000101:	sigmoid = 21'b000000101101011100000;
		14'b11011100000110:	sigmoid = 21'b000000101101100001101;
		14'b11011100000111:	sigmoid = 21'b000000101101100111010;
		14'b11011100001000:	sigmoid = 21'b000000101101101101000;
		14'b11011100001001:	sigmoid = 21'b000000101101110010101;
		14'b11011100001010:	sigmoid = 21'b000000101101111000010;
		14'b11011100001011:	sigmoid = 21'b000000101101111110000;
		14'b11011100001100:	sigmoid = 21'b000000101110000011101;
		14'b11011100001101:	sigmoid = 21'b000000101110001001011;
		14'b11011100001110:	sigmoid = 21'b000000101110001111000;
		14'b11011100001111:	sigmoid = 21'b000000101110010100110;
		14'b11011100010000:	sigmoid = 21'b000000101110011010100;
		14'b11011100010001:	sigmoid = 21'b000000101110100000010;
		14'b11011100010010:	sigmoid = 21'b000000101110100110000;
		14'b11011100010011:	sigmoid = 21'b000000101110101011110;
		14'b11011100010100:	sigmoid = 21'b000000101110110001100;
		14'b11011100010101:	sigmoid = 21'b000000101110110111010;
		14'b11011100010110:	sigmoid = 21'b000000101110111101001;
		14'b11011100010111:	sigmoid = 21'b000000101111000010111;
		14'b11011100011000:	sigmoid = 21'b000000101111001000110;
		14'b11011100011001:	sigmoid = 21'b000000101111001110100;
		14'b11011100011010:	sigmoid = 21'b000000101111010100011;
		14'b11011100011011:	sigmoid = 21'b000000101111011010010;
		14'b11011100011100:	sigmoid = 21'b000000101111100000001;
		14'b11011100011101:	sigmoid = 21'b000000101111100110000;
		14'b11011100011110:	sigmoid = 21'b000000101111101011111;
		14'b11011100011111:	sigmoid = 21'b000000101111110001110;
		14'b11011100100000:	sigmoid = 21'b000000101111110111101;
		14'b11011100100001:	sigmoid = 21'b000000101111111101101;
		14'b11011100100010:	sigmoid = 21'b000000110000000011100;
		14'b11011100100011:	sigmoid = 21'b000000110000001001100;
		14'b11011100100100:	sigmoid = 21'b000000110000001111011;
		14'b11011100100101:	sigmoid = 21'b000000110000010101011;
		14'b11011100100110:	sigmoid = 21'b000000110000011011011;
		14'b11011100100111:	sigmoid = 21'b000000110000100001011;
		14'b11011100101000:	sigmoid = 21'b000000110000100111011;
		14'b11011100101001:	sigmoid = 21'b000000110000101101011;
		14'b11011100101010:	sigmoid = 21'b000000110000110011011;
		14'b11011100101011:	sigmoid = 21'b000000110000111001011;
		14'b11011100101100:	sigmoid = 21'b000000110000111111100;
		14'b11011100101101:	sigmoid = 21'b000000110001000101100;
		14'b11011100101110:	sigmoid = 21'b000000110001001011101;
		14'b11011100101111:	sigmoid = 21'b000000110001010001101;
		14'b11011100110000:	sigmoid = 21'b000000110001010111110;
		14'b11011100110001:	sigmoid = 21'b000000110001011101111;
		14'b11011100110010:	sigmoid = 21'b000000110001100100000;
		14'b11011100110011:	sigmoid = 21'b000000110001101010001;
		14'b11011100110100:	sigmoid = 21'b000000110001110000010;
		14'b11011100110101:	sigmoid = 21'b000000110001110110011;
		14'b11011100110110:	sigmoid = 21'b000000110001111100100;
		14'b11011100110111:	sigmoid = 21'b000000110010000010110;
		14'b11011100111000:	sigmoid = 21'b000000110010001000111;
		14'b11011100111001:	sigmoid = 21'b000000110010001111001;
		14'b11011100111010:	sigmoid = 21'b000000110010010101011;
		14'b11011100111011:	sigmoid = 21'b000000110010011011100;
		14'b11011100111100:	sigmoid = 21'b000000110010100001110;
		14'b11011100111101:	sigmoid = 21'b000000110010101000000;
		14'b11011100111110:	sigmoid = 21'b000000110010101110010;
		14'b11011100111111:	sigmoid = 21'b000000110010110100100;
		14'b11011101000000:	sigmoid = 21'b000000110010111010111;
		14'b11011101000001:	sigmoid = 21'b000000110011000001001;
		14'b11011101000010:	sigmoid = 21'b000000110011000111011;
		14'b11011101000011:	sigmoid = 21'b000000110011001101110;
		14'b11011101000100:	sigmoid = 21'b000000110011010100000;
		14'b11011101000101:	sigmoid = 21'b000000110011011010011;
		14'b11011101000110:	sigmoid = 21'b000000110011100000110;
		14'b11011101000111:	sigmoid = 21'b000000110011100111001;
		14'b11011101001000:	sigmoid = 21'b000000110011101101100;
		14'b11011101001001:	sigmoid = 21'b000000110011110011111;
		14'b11011101001010:	sigmoid = 21'b000000110011111010010;
		14'b11011101001011:	sigmoid = 21'b000000110100000000110;
		14'b11011101001100:	sigmoid = 21'b000000110100000111001;
		14'b11011101001101:	sigmoid = 21'b000000110100001101100;
		14'b11011101001110:	sigmoid = 21'b000000110100010100000;
		14'b11011101001111:	sigmoid = 21'b000000110100011010100;
		14'b11011101010000:	sigmoid = 21'b000000110100100001000;
		14'b11011101010001:	sigmoid = 21'b000000110100100111011;
		14'b11011101010010:	sigmoid = 21'b000000110100101101111;
		14'b11011101010011:	sigmoid = 21'b000000110100110100100;
		14'b11011101010100:	sigmoid = 21'b000000110100111011000;
		14'b11011101010101:	sigmoid = 21'b000000110101000001100;
		14'b11011101010110:	sigmoid = 21'b000000110101001000000;
		14'b11011101010111:	sigmoid = 21'b000000110101001110101;
		14'b11011101011000:	sigmoid = 21'b000000110101010101001;
		14'b11011101011001:	sigmoid = 21'b000000110101011011110;
		14'b11011101011010:	sigmoid = 21'b000000110101100010011;
		14'b11011101011011:	sigmoid = 21'b000000110101101001000;
		14'b11011101011100:	sigmoid = 21'b000000110101101111101;
		14'b11011101011101:	sigmoid = 21'b000000110101110110010;
		14'b11011101011110:	sigmoid = 21'b000000110101111100111;
		14'b11011101011111:	sigmoid = 21'b000000110110000011100;
		14'b11011101100000:	sigmoid = 21'b000000110110001010010;
		14'b11011101100001:	sigmoid = 21'b000000110110010000111;
		14'b11011101100010:	sigmoid = 21'b000000110110010111101;
		14'b11011101100011:	sigmoid = 21'b000000110110011110011;
		14'b11011101100100:	sigmoid = 21'b000000110110100101000;
		14'b11011101100101:	sigmoid = 21'b000000110110101011110;
		14'b11011101100110:	sigmoid = 21'b000000110110110010100;
		14'b11011101100111:	sigmoid = 21'b000000110110111001010;
		14'b11011101101000:	sigmoid = 21'b000000110111000000001;
		14'b11011101101001:	sigmoid = 21'b000000110111000110111;
		14'b11011101101010:	sigmoid = 21'b000000110111001101101;
		14'b11011101101011:	sigmoid = 21'b000000110111010100100;
		14'b11011101101100:	sigmoid = 21'b000000110111011011010;
		14'b11011101101101:	sigmoid = 21'b000000110111100010001;
		14'b11011101101110:	sigmoid = 21'b000000110111101001000;
		14'b11011101101111:	sigmoid = 21'b000000110111101111111;
		14'b11011101110000:	sigmoid = 21'b000000110111110110110;
		14'b11011101110001:	sigmoid = 21'b000000110111111101101;
		14'b11011101110010:	sigmoid = 21'b000000111000000100100;
		14'b11011101110011:	sigmoid = 21'b000000111000001011100;
		14'b11011101110100:	sigmoid = 21'b000000111000010010011;
		14'b11011101110101:	sigmoid = 21'b000000111000011001011;
		14'b11011101110110:	sigmoid = 21'b000000111000100000010;
		14'b11011101110111:	sigmoid = 21'b000000111000100111010;
		14'b11011101111000:	sigmoid = 21'b000000111000101110010;
		14'b11011101111001:	sigmoid = 21'b000000111000110101010;
		14'b11011101111010:	sigmoid = 21'b000000111000111100010;
		14'b11011101111011:	sigmoid = 21'b000000111001000011010;
		14'b11011101111100:	sigmoid = 21'b000000111001001010011;
		14'b11011101111101:	sigmoid = 21'b000000111001010001011;
		14'b11011101111110:	sigmoid = 21'b000000111001011000100;
		14'b11011101111111:	sigmoid = 21'b000000111001011111100;
		14'b11011110000000:	sigmoid = 21'b000000111001100110101;
		14'b11011110000001:	sigmoid = 21'b000000111001101101110;
		14'b11011110000010:	sigmoid = 21'b000000111001110100111;
		14'b11011110000011:	sigmoid = 21'b000000111001111100000;
		14'b11011110000100:	sigmoid = 21'b000000111010000011001;
		14'b11011110000101:	sigmoid = 21'b000000111010001010010;
		14'b11011110000110:	sigmoid = 21'b000000111010010001100;
		14'b11011110000111:	sigmoid = 21'b000000111010011000101;
		14'b11011110001000:	sigmoid = 21'b000000111010011111111;
		14'b11011110001001:	sigmoid = 21'b000000111010100111001;
		14'b11011110001010:	sigmoid = 21'b000000111010101110010;
		14'b11011110001011:	sigmoid = 21'b000000111010110101100;
		14'b11011110001100:	sigmoid = 21'b000000111010111100110;
		14'b11011110001101:	sigmoid = 21'b000000111011000100001;
		14'b11011110001110:	sigmoid = 21'b000000111011001011011;
		14'b11011110001111:	sigmoid = 21'b000000111011010010101;
		14'b11011110010000:	sigmoid = 21'b000000111011011010000;
		14'b11011110010001:	sigmoid = 21'b000000111011100001010;
		14'b11011110010010:	sigmoid = 21'b000000111011101000101;
		14'b11011110010011:	sigmoid = 21'b000000111011110000000;
		14'b11011110010100:	sigmoid = 21'b000000111011110111011;
		14'b11011110010101:	sigmoid = 21'b000000111011111110110;
		14'b11011110010110:	sigmoid = 21'b000000111100000110001;
		14'b11011110010111:	sigmoid = 21'b000000111100001101100;
		14'b11011110011000:	sigmoid = 21'b000000111100010101000;
		14'b11011110011001:	sigmoid = 21'b000000111100011100011;
		14'b11011110011010:	sigmoid = 21'b000000111100100011111;
		14'b11011110011011:	sigmoid = 21'b000000111100101011010;
		14'b11011110011100:	sigmoid = 21'b000000111100110010110;
		14'b11011110011101:	sigmoid = 21'b000000111100111010010;
		14'b11011110011110:	sigmoid = 21'b000000111101000001110;
		14'b11011110011111:	sigmoid = 21'b000000111101001001010;
		14'b11011110100000:	sigmoid = 21'b000000111101010000111;
		14'b11011110100001:	sigmoid = 21'b000000111101011000011;
		14'b11011110100010:	sigmoid = 21'b000000111101100000000;
		14'b11011110100011:	sigmoid = 21'b000000111101100111100;
		14'b11011110100100:	sigmoid = 21'b000000111101101111001;
		14'b11011110100101:	sigmoid = 21'b000000111101110110110;
		14'b11011110100110:	sigmoid = 21'b000000111101111110011;
		14'b11011110100111:	sigmoid = 21'b000000111110000110000;
		14'b11011110101000:	sigmoid = 21'b000000111110001101101;
		14'b11011110101001:	sigmoid = 21'b000000111110010101011;
		14'b11011110101010:	sigmoid = 21'b000000111110011101000;
		14'b11011110101011:	sigmoid = 21'b000000111110100100110;
		14'b11011110101100:	sigmoid = 21'b000000111110101100011;
		14'b11011110101101:	sigmoid = 21'b000000111110110100001;
		14'b11011110101110:	sigmoid = 21'b000000111110111011111;
		14'b11011110101111:	sigmoid = 21'b000000111111000011101;
		14'b11011110110000:	sigmoid = 21'b000000111111001011011;
		14'b11011110110001:	sigmoid = 21'b000000111111010011001;
		14'b11011110110010:	sigmoid = 21'b000000111111011011000;
		14'b11011110110011:	sigmoid = 21'b000000111111100010110;
		14'b11011110110100:	sigmoid = 21'b000000111111101010101;
		14'b11011110110101:	sigmoid = 21'b000000111111110010100;
		14'b11011110110110:	sigmoid = 21'b000000111111111010010;
		14'b11011110110111:	sigmoid = 21'b000001000000000010001;
		14'b11011110111000:	sigmoid = 21'b000001000000001010001;
		14'b11011110111001:	sigmoid = 21'b000001000000010010000;
		14'b11011110111010:	sigmoid = 21'b000001000000011001111;
		14'b11011110111011:	sigmoid = 21'b000001000000100001111;
		14'b11011110111100:	sigmoid = 21'b000001000000101001110;
		14'b11011110111101:	sigmoid = 21'b000001000000110001110;
		14'b11011110111110:	sigmoid = 21'b000001000000111001110;
		14'b11011110111111:	sigmoid = 21'b000001000001000001110;
		14'b11011111000000:	sigmoid = 21'b000001000001001001110;
		14'b11011111000001:	sigmoid = 21'b000001000001010001110;
		14'b11011111000010:	sigmoid = 21'b000001000001011001110;
		14'b11011111000011:	sigmoid = 21'b000001000001100001111;
		14'b11011111000100:	sigmoid = 21'b000001000001101001111;
		14'b11011111000101:	sigmoid = 21'b000001000001110010000;
		14'b11011111000110:	sigmoid = 21'b000001000001111010001;
		14'b11011111000111:	sigmoid = 21'b000001000010000010001;
		14'b11011111001000:	sigmoid = 21'b000001000010001010010;
		14'b11011111001001:	sigmoid = 21'b000001000010010010100;
		14'b11011111001010:	sigmoid = 21'b000001000010011010101;
		14'b11011111001011:	sigmoid = 21'b000001000010100010110;
		14'b11011111001100:	sigmoid = 21'b000001000010101011000;
		14'b11011111001101:	sigmoid = 21'b000001000010110011001;
		14'b11011111001110:	sigmoid = 21'b000001000010111011011;
		14'b11011111001111:	sigmoid = 21'b000001000011000011101;
		14'b11011111010000:	sigmoid = 21'b000001000011001011111;
		14'b11011111010001:	sigmoid = 21'b000001000011010100001;
		14'b11011111010010:	sigmoid = 21'b000001000011011100100;
		14'b11011111010011:	sigmoid = 21'b000001000011100100110;
		14'b11011111010100:	sigmoid = 21'b000001000011101101000;
		14'b11011111010101:	sigmoid = 21'b000001000011110101011;
		14'b11011111010110:	sigmoid = 21'b000001000011111101110;
		14'b11011111010111:	sigmoid = 21'b000001000100000110001;
		14'b11011111011000:	sigmoid = 21'b000001000100001110100;
		14'b11011111011001:	sigmoid = 21'b000001000100010110111;
		14'b11011111011010:	sigmoid = 21'b000001000100011111010;
		14'b11011111011011:	sigmoid = 21'b000001000100100111110;
		14'b11011111011100:	sigmoid = 21'b000001000100110000001;
		14'b11011111011101:	sigmoid = 21'b000001000100111000101;
		14'b11011111011110:	sigmoid = 21'b000001000101000001001;
		14'b11011111011111:	sigmoid = 21'b000001000101001001101;
		14'b11011111100000:	sigmoid = 21'b000001000101010010001;
		14'b11011111100001:	sigmoid = 21'b000001000101011010101;
		14'b11011111100010:	sigmoid = 21'b000001000101100011001;
		14'b11011111100011:	sigmoid = 21'b000001000101101011110;
		14'b11011111100100:	sigmoid = 21'b000001000101110100010;
		14'b11011111100101:	sigmoid = 21'b000001000101111100111;
		14'b11011111100110:	sigmoid = 21'b000001000110000101100;
		14'b11011111100111:	sigmoid = 21'b000001000110001110001;
		14'b11011111101000:	sigmoid = 21'b000001000110010110110;
		14'b11011111101001:	sigmoid = 21'b000001000110011111011;
		14'b11011111101010:	sigmoid = 21'b000001000110101000000;
		14'b11011111101011:	sigmoid = 21'b000001000110110000110;
		14'b11011111101100:	sigmoid = 21'b000001000110111001011;
		14'b11011111101101:	sigmoid = 21'b000001000111000010001;
		14'b11011111101110:	sigmoid = 21'b000001000111001010111;
		14'b11011111101111:	sigmoid = 21'b000001000111010011101;
		14'b11011111110000:	sigmoid = 21'b000001000111011100011;
		14'b11011111110001:	sigmoid = 21'b000001000111100101001;
		14'b11011111110010:	sigmoid = 21'b000001000111101110000;
		14'b11011111110011:	sigmoid = 21'b000001000111110110110;
		14'b11011111110100:	sigmoid = 21'b000001000111111111101;
		14'b11011111110101:	sigmoid = 21'b000001001000001000100;
		14'b11011111110110:	sigmoid = 21'b000001001000010001011;
		14'b11011111110111:	sigmoid = 21'b000001001000011010010;
		14'b11011111111000:	sigmoid = 21'b000001001000100011001;
		14'b11011111111001:	sigmoid = 21'b000001001000101100000;
		14'b11011111111010:	sigmoid = 21'b000001001000110101000;
		14'b11011111111011:	sigmoid = 21'b000001001000111101111;
		14'b11011111111100:	sigmoid = 21'b000001001001000110111;
		14'b11011111111101:	sigmoid = 21'b000001001001001111111;
		14'b11011111111110:	sigmoid = 21'b000001001001011000111;
		14'b11011111111111:	sigmoid = 21'b000001001001100001111;
		14'b11100000000000:	sigmoid = 21'b000001001001101010111;
		14'b11100000000001:	sigmoid = 21'b000001001001110100000;
		14'b11100000000010:	sigmoid = 21'b000001001001111101000;
		14'b11100000000011:	sigmoid = 21'b000001001010000110001;
		14'b11100000000100:	sigmoid = 21'b000001001010001111010;
		14'b11100000000101:	sigmoid = 21'b000001001010011000011;
		14'b11100000000110:	sigmoid = 21'b000001001010100001100;
		14'b11100000000111:	sigmoid = 21'b000001001010101010101;
		14'b11100000001000:	sigmoid = 21'b000001001010110011110;
		14'b11100000001001:	sigmoid = 21'b000001001010111101000;
		14'b11100000001010:	sigmoid = 21'b000001001011000110010;
		14'b11100000001011:	sigmoid = 21'b000001001011001111011;
		14'b11100000001100:	sigmoid = 21'b000001001011011000101;
		14'b11100000001101:	sigmoid = 21'b000001001011100001111;
		14'b11100000001110:	sigmoid = 21'b000001001011101011010;
		14'b11100000001111:	sigmoid = 21'b000001001011110100100;
		14'b11100000010000:	sigmoid = 21'b000001001011111101110;
		14'b11100000010001:	sigmoid = 21'b000001001100000111001;
		14'b11100000010010:	sigmoid = 21'b000001001100010000100;
		14'b11100000010011:	sigmoid = 21'b000001001100011001111;
		14'b11100000010100:	sigmoid = 21'b000001001100100011010;
		14'b11100000010101:	sigmoid = 21'b000001001100101100101;
		14'b11100000010110:	sigmoid = 21'b000001001100110110000;
		14'b11100000010111:	sigmoid = 21'b000001001100111111100;
		14'b11100000011000:	sigmoid = 21'b000001001101001000111;
		14'b11100000011001:	sigmoid = 21'b000001001101010010011;
		14'b11100000011010:	sigmoid = 21'b000001001101011011111;
		14'b11100000011011:	sigmoid = 21'b000001001101100101011;
		14'b11100000011100:	sigmoid = 21'b000001001101101110111;
		14'b11100000011101:	sigmoid = 21'b000001001101111000100;
		14'b11100000011110:	sigmoid = 21'b000001001110000010000;
		14'b11100000011111:	sigmoid = 21'b000001001110001011101;
		14'b11100000100000:	sigmoid = 21'b000001001110010101010;
		14'b11100000100001:	sigmoid = 21'b000001001110011110110;
		14'b11100000100010:	sigmoid = 21'b000001001110101000011;
		14'b11100000100011:	sigmoid = 21'b000001001110110010001;
		14'b11100000100100:	sigmoid = 21'b000001001110111011110;
		14'b11100000100101:	sigmoid = 21'b000001001111000101011;
		14'b11100000100110:	sigmoid = 21'b000001001111001111001;
		14'b11100000100111:	sigmoid = 21'b000001001111011000111;
		14'b11100000101000:	sigmoid = 21'b000001001111100010101;
		14'b11100000101001:	sigmoid = 21'b000001001111101100011;
		14'b11100000101010:	sigmoid = 21'b000001001111110110001;
		14'b11100000101011:	sigmoid = 21'b000001001111111111111;
		14'b11100000101100:	sigmoid = 21'b000001010000001001110;
		14'b11100000101101:	sigmoid = 21'b000001010000010011101;
		14'b11100000101110:	sigmoid = 21'b000001010000011101011;
		14'b11100000101111:	sigmoid = 21'b000001010000100111010;
		14'b11100000110000:	sigmoid = 21'b000001010000110001010;
		14'b11100000110001:	sigmoid = 21'b000001010000111011001;
		14'b11100000110010:	sigmoid = 21'b000001010001000101000;
		14'b11100000110011:	sigmoid = 21'b000001010001001111000;
		14'b11100000110100:	sigmoid = 21'b000001010001011000111;
		14'b11100000110101:	sigmoid = 21'b000001010001100010111;
		14'b11100000110110:	sigmoid = 21'b000001010001101100111;
		14'b11100000110111:	sigmoid = 21'b000001010001110110111;
		14'b11100000111000:	sigmoid = 21'b000001010010000001000;
		14'b11100000111001:	sigmoid = 21'b000001010010001011000;
		14'b11100000111010:	sigmoid = 21'b000001010010010101001;
		14'b11100000111011:	sigmoid = 21'b000001010010011111010;
		14'b11100000111100:	sigmoid = 21'b000001010010101001010;
		14'b11100000111101:	sigmoid = 21'b000001010010110011011;
		14'b11100000111110:	sigmoid = 21'b000001010010111101101;
		14'b11100000111111:	sigmoid = 21'b000001010011000111110;
		14'b11100001000000:	sigmoid = 21'b000001010011010010000;
		14'b11100001000001:	sigmoid = 21'b000001010011011100001;
		14'b11100001000010:	sigmoid = 21'b000001010011100110011;
		14'b11100001000011:	sigmoid = 21'b000001010011110000101;
		14'b11100001000100:	sigmoid = 21'b000001010011111010111;
		14'b11100001000101:	sigmoid = 21'b000001010100000101001;
		14'b11100001000110:	sigmoid = 21'b000001010100001111100;
		14'b11100001000111:	sigmoid = 21'b000001010100011001110;
		14'b11100001001000:	sigmoid = 21'b000001010100100100001;
		14'b11100001001001:	sigmoid = 21'b000001010100101110100;
		14'b11100001001010:	sigmoid = 21'b000001010100111000111;
		14'b11100001001011:	sigmoid = 21'b000001010101000011010;
		14'b11100001001100:	sigmoid = 21'b000001010101001101110;
		14'b11100001001101:	sigmoid = 21'b000001010101011000001;
		14'b11100001001110:	sigmoid = 21'b000001010101100010101;
		14'b11100001001111:	sigmoid = 21'b000001010101101101001;
		14'b11100001010000:	sigmoid = 21'b000001010101110111101;
		14'b11100001010001:	sigmoid = 21'b000001010110000010001;
		14'b11100001010010:	sigmoid = 21'b000001010110001100101;
		14'b11100001010011:	sigmoid = 21'b000001010110010111010;
		14'b11100001010100:	sigmoid = 21'b000001010110100001110;
		14'b11100001010101:	sigmoid = 21'b000001010110101100011;
		14'b11100001010110:	sigmoid = 21'b000001010110110111000;
		14'b11100001010111:	sigmoid = 21'b000001010111000001101;
		14'b11100001011000:	sigmoid = 21'b000001010111001100010;
		14'b11100001011001:	sigmoid = 21'b000001010111010111000;
		14'b11100001011010:	sigmoid = 21'b000001010111100001101;
		14'b11100001011011:	sigmoid = 21'b000001010111101100011;
		14'b11100001011100:	sigmoid = 21'b000001010111110111001;
		14'b11100001011101:	sigmoid = 21'b000001011000000001111;
		14'b11100001011110:	sigmoid = 21'b000001011000001100101;
		14'b11100001011111:	sigmoid = 21'b000001011000010111100;
		14'b11100001100000:	sigmoid = 21'b000001011000100010010;
		14'b11100001100001:	sigmoid = 21'b000001011000101101001;
		14'b11100001100010:	sigmoid = 21'b000001011000111000000;
		14'b11100001100011:	sigmoid = 21'b000001011001000010111;
		14'b11100001100100:	sigmoid = 21'b000001011001001101110;
		14'b11100001100101:	sigmoid = 21'b000001011001011000101;
		14'b11100001100110:	sigmoid = 21'b000001011001100011101;
		14'b11100001100111:	sigmoid = 21'b000001011001101110100;
		14'b11100001101000:	sigmoid = 21'b000001011001111001100;
		14'b11100001101001:	sigmoid = 21'b000001011010000100100;
		14'b11100001101010:	sigmoid = 21'b000001011010001111101;
		14'b11100001101011:	sigmoid = 21'b000001011010011010101;
		14'b11100001101100:	sigmoid = 21'b000001011010100101101;
		14'b11100001101101:	sigmoid = 21'b000001011010110000110;
		14'b11100001101110:	sigmoid = 21'b000001011010111011111;
		14'b11100001101111:	sigmoid = 21'b000001011011000111000;
		14'b11100001110000:	sigmoid = 21'b000001011011010010001;
		14'b11100001110001:	sigmoid = 21'b000001011011011101010;
		14'b11100001110010:	sigmoid = 21'b000001011011101000100;
		14'b11100001110011:	sigmoid = 21'b000001011011110011110;
		14'b11100001110100:	sigmoid = 21'b000001011011111110111;
		14'b11100001110101:	sigmoid = 21'b000001011100001010001;
		14'b11100001110110:	sigmoid = 21'b000001011100010101100;
		14'b11100001110111:	sigmoid = 21'b000001011100100000110;
		14'b11100001111000:	sigmoid = 21'b000001011100101100000;
		14'b11100001111001:	sigmoid = 21'b000001011100110111011;
		14'b11100001111010:	sigmoid = 21'b000001011101000010110;
		14'b11100001111011:	sigmoid = 21'b000001011101001110001;
		14'b11100001111100:	sigmoid = 21'b000001011101011001100;
		14'b11100001111101:	sigmoid = 21'b000001011101100100111;
		14'b11100001111110:	sigmoid = 21'b000001011101110000011;
		14'b11100001111111:	sigmoid = 21'b000001011101111011111;
		14'b11100010000000:	sigmoid = 21'b000001011110000111011;
		14'b11100010000001:	sigmoid = 21'b000001011110010010111;
		14'b11100010000010:	sigmoid = 21'b000001011110011110011;
		14'b11100010000011:	sigmoid = 21'b000001011110101001111;
		14'b11100010000100:	sigmoid = 21'b000001011110110101100;
		14'b11100010000101:	sigmoid = 21'b000001011111000001000;
		14'b11100010000110:	sigmoid = 21'b000001011111001100101;
		14'b11100010000111:	sigmoid = 21'b000001011111011000010;
		14'b11100010001000:	sigmoid = 21'b000001011111100100000;
		14'b11100010001001:	sigmoid = 21'b000001011111101111101;
		14'b11100010001010:	sigmoid = 21'b000001011111111011011;
		14'b11100010001011:	sigmoid = 21'b000001100000000111000;
		14'b11100010001100:	sigmoid = 21'b000001100000010010110;
		14'b11100010001101:	sigmoid = 21'b000001100000011110101;
		14'b11100010001110:	sigmoid = 21'b000001100000101010011;
		14'b11100010001111:	sigmoid = 21'b000001100000110110001;
		14'b11100010010000:	sigmoid = 21'b000001100001000010000;
		14'b11100010010001:	sigmoid = 21'b000001100001001101111;
		14'b11100010010010:	sigmoid = 21'b000001100001011001110;
		14'b11100010010011:	sigmoid = 21'b000001100001100101101;
		14'b11100010010100:	sigmoid = 21'b000001100001110001100;
		14'b11100010010101:	sigmoid = 21'b000001100001111101100;
		14'b11100010010110:	sigmoid = 21'b000001100010001001100;
		14'b11100010010111:	sigmoid = 21'b000001100010010101011;
		14'b11100010011000:	sigmoid = 21'b000001100010100001011;
		14'b11100010011001:	sigmoid = 21'b000001100010101101100;
		14'b11100010011010:	sigmoid = 21'b000001100010111001100;
		14'b11100010011011:	sigmoid = 21'b000001100011000101101;
		14'b11100010011100:	sigmoid = 21'b000001100011010001110;
		14'b11100010011101:	sigmoid = 21'b000001100011011101110;
		14'b11100010011110:	sigmoid = 21'b000001100011101010000;
		14'b11100010011111:	sigmoid = 21'b000001100011110110001;
		14'b11100010100000:	sigmoid = 21'b000001100100000010010;
		14'b11100010100001:	sigmoid = 21'b000001100100001110100;
		14'b11100010100010:	sigmoid = 21'b000001100100011010110;
		14'b11100010100011:	sigmoid = 21'b000001100100100111000;
		14'b11100010100100:	sigmoid = 21'b000001100100110011010;
		14'b11100010100101:	sigmoid = 21'b000001100100111111101;
		14'b11100010100110:	sigmoid = 21'b000001100101001011111;
		14'b11100010100111:	sigmoid = 21'b000001100101011000010;
		14'b11100010101000:	sigmoid = 21'b000001100101100100101;
		14'b11100010101001:	sigmoid = 21'b000001100101110001000;
		14'b11100010101010:	sigmoid = 21'b000001100101111101011;
		14'b11100010101011:	sigmoid = 21'b000001100110001001111;
		14'b11100010101100:	sigmoid = 21'b000001100110010110011;
		14'b11100010101101:	sigmoid = 21'b000001100110100010111;
		14'b11100010101110:	sigmoid = 21'b000001100110101111011;
		14'b11100010101111:	sigmoid = 21'b000001100110111011111;
		14'b11100010110000:	sigmoid = 21'b000001100111001000011;
		14'b11100010110001:	sigmoid = 21'b000001100111010101000;
		14'b11100010110010:	sigmoid = 21'b000001100111100001101;
		14'b11100010110011:	sigmoid = 21'b000001100111101110010;
		14'b11100010110100:	sigmoid = 21'b000001100111111010111;
		14'b11100010110101:	sigmoid = 21'b000001101000000111100;
		14'b11100010110110:	sigmoid = 21'b000001101000010100010;
		14'b11100010110111:	sigmoid = 21'b000001101000100001000;
		14'b11100010111000:	sigmoid = 21'b000001101000101101110;
		14'b11100010111001:	sigmoid = 21'b000001101000111010100;
		14'b11100010111010:	sigmoid = 21'b000001101001000111010;
		14'b11100010111011:	sigmoid = 21'b000001101001010100001;
		14'b11100010111100:	sigmoid = 21'b000001101001100000111;
		14'b11100010111101:	sigmoid = 21'b000001101001101101110;
		14'b11100010111110:	sigmoid = 21'b000001101001111010101;
		14'b11100010111111:	sigmoid = 21'b000001101010000111101;
		14'b11100011000000:	sigmoid = 21'b000001101010010100100;
		14'b11100011000001:	sigmoid = 21'b000001101010100001100;
		14'b11100011000010:	sigmoid = 21'b000001101010101110100;
		14'b11100011000011:	sigmoid = 21'b000001101010111011100;
		14'b11100011000100:	sigmoid = 21'b000001101011001000100;
		14'b11100011000101:	sigmoid = 21'b000001101011010101100;
		14'b11100011000110:	sigmoid = 21'b000001101011100010101;
		14'b11100011000111:	sigmoid = 21'b000001101011101111110;
		14'b11100011001000:	sigmoid = 21'b000001101011111100111;
		14'b11100011001001:	sigmoid = 21'b000001101100001010000;
		14'b11100011001010:	sigmoid = 21'b000001101100010111001;
		14'b11100011001011:	sigmoid = 21'b000001101100100100011;
		14'b11100011001100:	sigmoid = 21'b000001101100110001101;
		14'b11100011001101:	sigmoid = 21'b000001101100111110111;
		14'b11100011001110:	sigmoid = 21'b000001101101001100001;
		14'b11100011001111:	sigmoid = 21'b000001101101011001011;
		14'b11100011010000:	sigmoid = 21'b000001101101100110110;
		14'b11100011010001:	sigmoid = 21'b000001101101110100001;
		14'b11100011010010:	sigmoid = 21'b000001101110000001100;
		14'b11100011010011:	sigmoid = 21'b000001101110001110111;
		14'b11100011010100:	sigmoid = 21'b000001101110011100010;
		14'b11100011010101:	sigmoid = 21'b000001101110101001110;
		14'b11100011010110:	sigmoid = 21'b000001101110110111001;
		14'b11100011010111:	sigmoid = 21'b000001101111000100101;
		14'b11100011011000:	sigmoid = 21'b000001101111010010010;
		14'b11100011011001:	sigmoid = 21'b000001101111011111110;
		14'b11100011011010:	sigmoid = 21'b000001101111101101010;
		14'b11100011011011:	sigmoid = 21'b000001101111111010111;
		14'b11100011011100:	sigmoid = 21'b000001110000001000100;
		14'b11100011011101:	sigmoid = 21'b000001110000010110001;
		14'b11100011011110:	sigmoid = 21'b000001110000100011111;
		14'b11100011011111:	sigmoid = 21'b000001110000110001100;
		14'b11100011100000:	sigmoid = 21'b000001110000111111010;
		14'b11100011100001:	sigmoid = 21'b000001110001001101000;
		14'b11100011100010:	sigmoid = 21'b000001110001011010110;
		14'b11100011100011:	sigmoid = 21'b000001110001101000101;
		14'b11100011100100:	sigmoid = 21'b000001110001110110011;
		14'b11100011100101:	sigmoid = 21'b000001110010000100010;
		14'b11100011100110:	sigmoid = 21'b000001110010010010001;
		14'b11100011100111:	sigmoid = 21'b000001110010100000000;
		14'b11100011101000:	sigmoid = 21'b000001110010101110000;
		14'b11100011101001:	sigmoid = 21'b000001110010111011111;
		14'b11100011101010:	sigmoid = 21'b000001110011001001111;
		14'b11100011101011:	sigmoid = 21'b000001110011010111111;
		14'b11100011101100:	sigmoid = 21'b000001110011100101111;
		14'b11100011101101:	sigmoid = 21'b000001110011110100000;
		14'b11100011101110:	sigmoid = 21'b000001110100000010000;
		14'b11100011101111:	sigmoid = 21'b000001110100010000001;
		14'b11100011110000:	sigmoid = 21'b000001110100011110010;
		14'b11100011110001:	sigmoid = 21'b000001110100101100011;
		14'b11100011110010:	sigmoid = 21'b000001110100111010101;
		14'b11100011110011:	sigmoid = 21'b000001110101001000111;
		14'b11100011110100:	sigmoid = 21'b000001110101010111001;
		14'b11100011110101:	sigmoid = 21'b000001110101100101011;
		14'b11100011110110:	sigmoid = 21'b000001110101110011101;
		14'b11100011110111:	sigmoid = 21'b000001110110000001111;
		14'b11100011111000:	sigmoid = 21'b000001110110010000010;
		14'b11100011111001:	sigmoid = 21'b000001110110011110101;
		14'b11100011111010:	sigmoid = 21'b000001110110101101000;
		14'b11100011111011:	sigmoid = 21'b000001110110111011100;
		14'b11100011111100:	sigmoid = 21'b000001110111001001111;
		14'b11100011111101:	sigmoid = 21'b000001110111011000011;
		14'b11100011111110:	sigmoid = 21'b000001110111100110111;
		14'b11100011111111:	sigmoid = 21'b000001110111110101011;
		14'b11100100000000:	sigmoid = 21'b000001111000000100000;
		14'b11100100000001:	sigmoid = 21'b000001111000010010100;
		14'b11100100000010:	sigmoid = 21'b000001111000100001001;
		14'b11100100000011:	sigmoid = 21'b000001111000101111110;
		14'b11100100000100:	sigmoid = 21'b000001111000111110100;
		14'b11100100000101:	sigmoid = 21'b000001111001001101001;
		14'b11100100000110:	sigmoid = 21'b000001111001011011111;
		14'b11100100000111:	sigmoid = 21'b000001111001101010101;
		14'b11100100001000:	sigmoid = 21'b000001111001111001011;
		14'b11100100001001:	sigmoid = 21'b000001111010001000001;
		14'b11100100001010:	sigmoid = 21'b000001111010010111000;
		14'b11100100001011:	sigmoid = 21'b000001111010100101111;
		14'b11100100001100:	sigmoid = 21'b000001111010110100110;
		14'b11100100001101:	sigmoid = 21'b000001111011000011101;
		14'b11100100001110:	sigmoid = 21'b000001111011010010100;
		14'b11100100001111:	sigmoid = 21'b000001111011100001100;
		14'b11100100010000:	sigmoid = 21'b000001111011110000100;
		14'b11100100010001:	sigmoid = 21'b000001111011111111100;
		14'b11100100010010:	sigmoid = 21'b000001111100001110101;
		14'b11100100010011:	sigmoid = 21'b000001111100011101101;
		14'b11100100010100:	sigmoid = 21'b000001111100101100110;
		14'b11100100010101:	sigmoid = 21'b000001111100111011111;
		14'b11100100010110:	sigmoid = 21'b000001111101001011000;
		14'b11100100010111:	sigmoid = 21'b000001111101011010010;
		14'b11100100011000:	sigmoid = 21'b000001111101101001011;
		14'b11100100011001:	sigmoid = 21'b000001111101111000101;
		14'b11100100011010:	sigmoid = 21'b000001111110000111111;
		14'b11100100011011:	sigmoid = 21'b000001111110010111010;
		14'b11100100011100:	sigmoid = 21'b000001111110100110100;
		14'b11100100011101:	sigmoid = 21'b000001111110110101111;
		14'b11100100011110:	sigmoid = 21'b000001111111000101010;
		14'b11100100011111:	sigmoid = 21'b000001111111010100101;
		14'b11100100100000:	sigmoid = 21'b000001111111100100001;
		14'b11100100100001:	sigmoid = 21'b000001111111110011101;
		14'b11100100100010:	sigmoid = 21'b000010000000000011000;
		14'b11100100100011:	sigmoid = 21'b000010000000010010101;
		14'b11100100100100:	sigmoid = 21'b000010000000100010001;
		14'b11100100100101:	sigmoid = 21'b000010000000110001110;
		14'b11100100100110:	sigmoid = 21'b000010000001000001010;
		14'b11100100100111:	sigmoid = 21'b000010000001010001000;
		14'b11100100101000:	sigmoid = 21'b000010000001100000101;
		14'b11100100101001:	sigmoid = 21'b000010000001110000010;
		14'b11100100101010:	sigmoid = 21'b000010000010000000000;
		14'b11100100101011:	sigmoid = 21'b000010000010001111110;
		14'b11100100101100:	sigmoid = 21'b000010000010011111100;
		14'b11100100101101:	sigmoid = 21'b000010000010101111011;
		14'b11100100101110:	sigmoid = 21'b000010000010111111001;
		14'b11100100101111:	sigmoid = 21'b000010000011001111000;
		14'b11100100110000:	sigmoid = 21'b000010000011011111000;
		14'b11100100110001:	sigmoid = 21'b000010000011101110111;
		14'b11100100110010:	sigmoid = 21'b000010000011111110111;
		14'b11100100110011:	sigmoid = 21'b000010000100001110110;
		14'b11100100110100:	sigmoid = 21'b000010000100011110110;
		14'b11100100110101:	sigmoid = 21'b000010000100101110111;
		14'b11100100110110:	sigmoid = 21'b000010000100111110111;
		14'b11100100110111:	sigmoid = 21'b000010000101001111000;
		14'b11100100111000:	sigmoid = 21'b000010000101011111001;
		14'b11100100111001:	sigmoid = 21'b000010000101101111010;
		14'b11100100111010:	sigmoid = 21'b000010000101111111100;
		14'b11100100111011:	sigmoid = 21'b000010000110001111110;
		14'b11100100111100:	sigmoid = 21'b000010000110100000000;
		14'b11100100111101:	sigmoid = 21'b000010000110110000010;
		14'b11100100111110:	sigmoid = 21'b000010000111000000100;
		14'b11100100111111:	sigmoid = 21'b000010000111010000111;
		14'b11100101000000:	sigmoid = 21'b000010000111100001010;
		14'b11100101000001:	sigmoid = 21'b000010000111110001101;
		14'b11100101000010:	sigmoid = 21'b000010001000000010000;
		14'b11100101000011:	sigmoid = 21'b000010001000010010100;
		14'b11100101000100:	sigmoid = 21'b000010001000100011000;
		14'b11100101000101:	sigmoid = 21'b000010001000110011100;
		14'b11100101000110:	sigmoid = 21'b000010001001000100000;
		14'b11100101000111:	sigmoid = 21'b000010001001010100101;
		14'b11100101001000:	sigmoid = 21'b000010001001100101010;
		14'b11100101001001:	sigmoid = 21'b000010001001110101111;
		14'b11100101001010:	sigmoid = 21'b000010001010000110100;
		14'b11100101001011:	sigmoid = 21'b000010001010010111010;
		14'b11100101001100:	sigmoid = 21'b000010001010101000000;
		14'b11100101001101:	sigmoid = 21'b000010001010111000110;
		14'b11100101001110:	sigmoid = 21'b000010001011001001100;
		14'b11100101001111:	sigmoid = 21'b000010001011011010010;
		14'b11100101010000:	sigmoid = 21'b000010001011101011001;
		14'b11100101010001:	sigmoid = 21'b000010001011111100000;
		14'b11100101010010:	sigmoid = 21'b000010001100001101000;
		14'b11100101010011:	sigmoid = 21'b000010001100011101111;
		14'b11100101010100:	sigmoid = 21'b000010001100101110111;
		14'b11100101010101:	sigmoid = 21'b000010001100111111111;
		14'b11100101010110:	sigmoid = 21'b000010001101010000111;
		14'b11100101010111:	sigmoid = 21'b000010001101100010000;
		14'b11100101011000:	sigmoid = 21'b000010001101110011000;
		14'b11100101011001:	sigmoid = 21'b000010001110000100001;
		14'b11100101011010:	sigmoid = 21'b000010001110010101011;
		14'b11100101011011:	sigmoid = 21'b000010001110100110100;
		14'b11100101011100:	sigmoid = 21'b000010001110110111110;
		14'b11100101011101:	sigmoid = 21'b000010001111001001000;
		14'b11100101011110:	sigmoid = 21'b000010001111011010010;
		14'b11100101011111:	sigmoid = 21'b000010001111101011101;
		14'b11100101100000:	sigmoid = 21'b000010001111111101000;
		14'b11100101100001:	sigmoid = 21'b000010010000001110011;
		14'b11100101100010:	sigmoid = 21'b000010010000011111110;
		14'b11100101100011:	sigmoid = 21'b000010010000110001001;
		14'b11100101100100:	sigmoid = 21'b000010010001000010101;
		14'b11100101100101:	sigmoid = 21'b000010010001010100001;
		14'b11100101100110:	sigmoid = 21'b000010010001100101110;
		14'b11100101100111:	sigmoid = 21'b000010010001110111010;
		14'b11100101101000:	sigmoid = 21'b000010010010001000111;
		14'b11100101101001:	sigmoid = 21'b000010010010011010100;
		14'b11100101101010:	sigmoid = 21'b000010010010101100001;
		14'b11100101101011:	sigmoid = 21'b000010010010111101111;
		14'b11100101101100:	sigmoid = 21'b000010010011001111101;
		14'b11100101101101:	sigmoid = 21'b000010010011100001011;
		14'b11100101101110:	sigmoid = 21'b000010010011110011001;
		14'b11100101101111:	sigmoid = 21'b000010010100000101000;
		14'b11100101110000:	sigmoid = 21'b000010010100010110110;
		14'b11100101110001:	sigmoid = 21'b000010010100101000110;
		14'b11100101110010:	sigmoid = 21'b000010010100111010101;
		14'b11100101110011:	sigmoid = 21'b000010010101001100101;
		14'b11100101110100:	sigmoid = 21'b000010010101011110100;
		14'b11100101110101:	sigmoid = 21'b000010010101110000101;
		14'b11100101110110:	sigmoid = 21'b000010010110000010101;
		14'b11100101110111:	sigmoid = 21'b000010010110010100110;
		14'b11100101111000:	sigmoid = 21'b000010010110100110111;
		14'b11100101111001:	sigmoid = 21'b000010010110111001000;
		14'b11100101111010:	sigmoid = 21'b000010010111001011001;
		14'b11100101111011:	sigmoid = 21'b000010010111011101011;
		14'b11100101111100:	sigmoid = 21'b000010010111101111101;
		14'b11100101111101:	sigmoid = 21'b000010011000000001111;
		14'b11100101111110:	sigmoid = 21'b000010011000010100010;
		14'b11100101111111:	sigmoid = 21'b000010011000100110101;
		14'b11100110000000:	sigmoid = 21'b000010011000111001000;
		14'b11100110000001:	sigmoid = 21'b000010011001001011011;
		14'b11100110000010:	sigmoid = 21'b000010011001011101111;
		14'b11100110000011:	sigmoid = 21'b000010011001110000010;
		14'b11100110000100:	sigmoid = 21'b000010011010000010111;
		14'b11100110000101:	sigmoid = 21'b000010011010010101011;
		14'b11100110000110:	sigmoid = 21'b000010011010101000000;
		14'b11100110000111:	sigmoid = 21'b000010011010111010100;
		14'b11100110001000:	sigmoid = 21'b000010011011001101010;
		14'b11100110001001:	sigmoid = 21'b000010011011011111111;
		14'b11100110001010:	sigmoid = 21'b000010011011110010101;
		14'b11100110001011:	sigmoid = 21'b000010011100000101011;
		14'b11100110001100:	sigmoid = 21'b000010011100011000001;
		14'b11100110001101:	sigmoid = 21'b000010011100101011000;
		14'b11100110001110:	sigmoid = 21'b000010011100111101111;
		14'b11100110001111:	sigmoid = 21'b000010011101010000110;
		14'b11100110010000:	sigmoid = 21'b000010011101100011101;
		14'b11100110010001:	sigmoid = 21'b000010011101110110101;
		14'b11100110010010:	sigmoid = 21'b000010011110001001100;
		14'b11100110010011:	sigmoid = 21'b000010011110011100101;
		14'b11100110010100:	sigmoid = 21'b000010011110101111101;
		14'b11100110010101:	sigmoid = 21'b000010011111000010110;
		14'b11100110010110:	sigmoid = 21'b000010011111010101111;
		14'b11100110010111:	sigmoid = 21'b000010011111101001000;
		14'b11100110011000:	sigmoid = 21'b000010011111111100010;
		14'b11100110011001:	sigmoid = 21'b000010100000001111100;
		14'b11100110011010:	sigmoid = 21'b000010100000100010110;
		14'b11100110011011:	sigmoid = 21'b000010100000110110000;
		14'b11100110011100:	sigmoid = 21'b000010100001001001011;
		14'b11100110011101:	sigmoid = 21'b000010100001011100110;
		14'b11100110011110:	sigmoid = 21'b000010100001110000001;
		14'b11100110011111:	sigmoid = 21'b000010100010000011100;
		14'b11100110100000:	sigmoid = 21'b000010100010010111000;
		14'b11100110100001:	sigmoid = 21'b000010100010101010100;
		14'b11100110100010:	sigmoid = 21'b000010100010111110001;
		14'b11100110100011:	sigmoid = 21'b000010100011010001101;
		14'b11100110100100:	sigmoid = 21'b000010100011100101010;
		14'b11100110100101:	sigmoid = 21'b000010100011111000111;
		14'b11100110100110:	sigmoid = 21'b000010100100001100101;
		14'b11100110100111:	sigmoid = 21'b000010100100100000011;
		14'b11100110101000:	sigmoid = 21'b000010100100110100001;
		14'b11100110101001:	sigmoid = 21'b000010100101000111111;
		14'b11100110101010:	sigmoid = 21'b000010100101011011110;
		14'b11100110101011:	sigmoid = 21'b000010100101101111100;
		14'b11100110101100:	sigmoid = 21'b000010100110000011100;
		14'b11100110101101:	sigmoid = 21'b000010100110010111011;
		14'b11100110101110:	sigmoid = 21'b000010100110101011011;
		14'b11100110101111:	sigmoid = 21'b000010100110111111011;
		14'b11100110110000:	sigmoid = 21'b000010100111010011011;
		14'b11100110110001:	sigmoid = 21'b000010100111100111100;
		14'b11100110110010:	sigmoid = 21'b000010100111111011101;
		14'b11100110110011:	sigmoid = 21'b000010101000001111110;
		14'b11100110110100:	sigmoid = 21'b000010101000100011111;
		14'b11100110110101:	sigmoid = 21'b000010101000111000001;
		14'b11100110110110:	sigmoid = 21'b000010101001001100011;
		14'b11100110110111:	sigmoid = 21'b000010101001100000110;
		14'b11100110111000:	sigmoid = 21'b000010101001110101000;
		14'b11100110111001:	sigmoid = 21'b000010101010001001011;
		14'b11100110111010:	sigmoid = 21'b000010101010011101110;
		14'b11100110111011:	sigmoid = 21'b000010101010110010010;
		14'b11100110111100:	sigmoid = 21'b000010101011000110110;
		14'b11100110111101:	sigmoid = 21'b000010101011011011010;
		14'b11100110111110:	sigmoid = 21'b000010101011101111110;
		14'b11100110111111:	sigmoid = 21'b000010101100000100011;
		14'b11100111000000:	sigmoid = 21'b000010101100011001000;
		14'b11100111000001:	sigmoid = 21'b000010101100101101101;
		14'b11100111000010:	sigmoid = 21'b000010101101000010011;
		14'b11100111000011:	sigmoid = 21'b000010101101010111001;
		14'b11100111000100:	sigmoid = 21'b000010101101101011111;
		14'b11100111000101:	sigmoid = 21'b000010101110000000101;
		14'b11100111000110:	sigmoid = 21'b000010101110010101100;
		14'b11100111000111:	sigmoid = 21'b000010101110101010011;
		14'b11100111001000:	sigmoid = 21'b000010101110111111010;
		14'b11100111001001:	sigmoid = 21'b000010101111010100010;
		14'b11100111001010:	sigmoid = 21'b000010101111101001010;
		14'b11100111001011:	sigmoid = 21'b000010101111111110010;
		14'b11100111001100:	sigmoid = 21'b000010110000010011011;
		14'b11100111001101:	sigmoid = 21'b000010110000101000100;
		14'b11100111001110:	sigmoid = 21'b000010110000111101101;
		14'b11100111001111:	sigmoid = 21'b000010110001010010110;
		14'b11100111010000:	sigmoid = 21'b000010110001101000000;
		14'b11100111010001:	sigmoid = 21'b000010110001111101010;
		14'b11100111010010:	sigmoid = 21'b000010110010010010101;
		14'b11100111010011:	sigmoid = 21'b000010110010100111111;
		14'b11100111010100:	sigmoid = 21'b000010110010111101010;
		14'b11100111010101:	sigmoid = 21'b000010110011010010110;
		14'b11100111010110:	sigmoid = 21'b000010110011101000001;
		14'b11100111010111:	sigmoid = 21'b000010110011111101101;
		14'b11100111011000:	sigmoid = 21'b000010110100010011001;
		14'b11100111011001:	sigmoid = 21'b000010110100101000110;
		14'b11100111011010:	sigmoid = 21'b000010110100111110011;
		14'b11100111011011:	sigmoid = 21'b000010110101010100000;
		14'b11100111011100:	sigmoid = 21'b000010110101101001101;
		14'b11100111011101:	sigmoid = 21'b000010110101111111011;
		14'b11100111011110:	sigmoid = 21'b000010110110010101001;
		14'b11100111011111:	sigmoid = 21'b000010110110101010111;
		14'b11100111100000:	sigmoid = 21'b000010110111000000110;
		14'b11100111100001:	sigmoid = 21'b000010110111010110101;
		14'b11100111100010:	sigmoid = 21'b000010110111101100100;
		14'b11100111100011:	sigmoid = 21'b000010111000000010100;
		14'b11100111100100:	sigmoid = 21'b000010111000011000100;
		14'b11100111100101:	sigmoid = 21'b000010111000101110100;
		14'b11100111100110:	sigmoid = 21'b000010111001000100101;
		14'b11100111100111:	sigmoid = 21'b000010111001011010110;
		14'b11100111101000:	sigmoid = 21'b000010111001110000111;
		14'b11100111101001:	sigmoid = 21'b000010111010000111000;
		14'b11100111101010:	sigmoid = 21'b000010111010011101010;
		14'b11100111101011:	sigmoid = 21'b000010111010110011100;
		14'b11100111101100:	sigmoid = 21'b000010111011001001111;
		14'b11100111101101:	sigmoid = 21'b000010111011100000001;
		14'b11100111101110:	sigmoid = 21'b000010111011110110100;
		14'b11100111101111:	sigmoid = 21'b000010111100001101000;
		14'b11100111110000:	sigmoid = 21'b000010111100100011100;
		14'b11100111110001:	sigmoid = 21'b000010111100111010000;
		14'b11100111110010:	sigmoid = 21'b000010111101010000100;
		14'b11100111110011:	sigmoid = 21'b000010111101100111001;
		14'b11100111110100:	sigmoid = 21'b000010111101111101110;
		14'b11100111110101:	sigmoid = 21'b000010111110010100011;
		14'b11100111110110:	sigmoid = 21'b000010111110101011001;
		14'b11100111110111:	sigmoid = 21'b000010111111000001111;
		14'b11100111111000:	sigmoid = 21'b000010111111011000101;
		14'b11100111111001:	sigmoid = 21'b000010111111101111011;
		14'b11100111111010:	sigmoid = 21'b000011000000000110010;
		14'b11100111111011:	sigmoid = 21'b000011000000011101010;
		14'b11100111111100:	sigmoid = 21'b000011000000110100001;
		14'b11100111111101:	sigmoid = 21'b000011000001001011001;
		14'b11100111111110:	sigmoid = 21'b000011000001100010001;
		14'b11100111111111:	sigmoid = 21'b000011000001111001010;
		14'b11101000000000:	sigmoid = 21'b000011000010010000011;
		14'b11101000000001:	sigmoid = 21'b000011000010100111100;
		14'b11101000000010:	sigmoid = 21'b000011000010111110110;
		14'b11101000000011:	sigmoid = 21'b000011000011010101111;
		14'b11101000000100:	sigmoid = 21'b000011000011101101010;
		14'b11101000000101:	sigmoid = 21'b000011000100000100100;
		14'b11101000000110:	sigmoid = 21'b000011000100011011111;
		14'b11101000000111:	sigmoid = 21'b000011000100110011010;
		14'b11101000001000:	sigmoid = 21'b000011000101001010110;
		14'b11101000001001:	sigmoid = 21'b000011000101100010001;
		14'b11101000001010:	sigmoid = 21'b000011000101111001110;
		14'b11101000001011:	sigmoid = 21'b000011000110010001010;
		14'b11101000001100:	sigmoid = 21'b000011000110101000111;
		14'b11101000001101:	sigmoid = 21'b000011000111000000100;
		14'b11101000001110:	sigmoid = 21'b000011000111011000010;
		14'b11101000001111:	sigmoid = 21'b000011000111110000000;
		14'b11101000010000:	sigmoid = 21'b000011001000000111110;
		14'b11101000010001:	sigmoid = 21'b000011001000011111100;
		14'b11101000010010:	sigmoid = 21'b000011001000110111011;
		14'b11101000010011:	sigmoid = 21'b000011001001001111010;
		14'b11101000010100:	sigmoid = 21'b000011001001100111010;
		14'b11101000010101:	sigmoid = 21'b000011001001111111010;
		14'b11101000010110:	sigmoid = 21'b000011001010010111010;
		14'b11101000010111:	sigmoid = 21'b000011001010101111010;
		14'b11101000011000:	sigmoid = 21'b000011001011000111011;
		14'b11101000011001:	sigmoid = 21'b000011001011011111100;
		14'b11101000011010:	sigmoid = 21'b000011001011110111110;
		14'b11101000011011:	sigmoid = 21'b000011001100010000000;
		14'b11101000011100:	sigmoid = 21'b000011001100101000010;
		14'b11101000011101:	sigmoid = 21'b000011001101000000101;
		14'b11101000011110:	sigmoid = 21'b000011001101011001000;
		14'b11101000011111:	sigmoid = 21'b000011001101110001011;
		14'b11101000100000:	sigmoid = 21'b000011001110001001110;
		14'b11101000100001:	sigmoid = 21'b000011001110100010010;
		14'b11101000100010:	sigmoid = 21'b000011001110111010111;
		14'b11101000100011:	sigmoid = 21'b000011001111010011011;
		14'b11101000100100:	sigmoid = 21'b000011001111101100000;
		14'b11101000100101:	sigmoid = 21'b000011010000000100110;
		14'b11101000100110:	sigmoid = 21'b000011010000011101011;
		14'b11101000100111:	sigmoid = 21'b000011010000110110001;
		14'b11101000101000:	sigmoid = 21'b000011010001001111000;
		14'b11101000101001:	sigmoid = 21'b000011010001100111110;
		14'b11101000101010:	sigmoid = 21'b000011010010000000110;
		14'b11101000101011:	sigmoid = 21'b000011010010011001101;
		14'b11101000101100:	sigmoid = 21'b000011010010110010101;
		14'b11101000101101:	sigmoid = 21'b000011010011001011101;
		14'b11101000101110:	sigmoid = 21'b000011010011100100101;
		14'b11101000101111:	sigmoid = 21'b000011010011111101110;
		14'b11101000110000:	sigmoid = 21'b000011010100010110111;
		14'b11101000110001:	sigmoid = 21'b000011010100110000001;
		14'b11101000110010:	sigmoid = 21'b000011010101001001011;
		14'b11101000110011:	sigmoid = 21'b000011010101100010101;
		14'b11101000110100:	sigmoid = 21'b000011010101111100000;
		14'b11101000110101:	sigmoid = 21'b000011010110010101010;
		14'b11101000110110:	sigmoid = 21'b000011010110101110110;
		14'b11101000110111:	sigmoid = 21'b000011010111001000001;
		14'b11101000111000:	sigmoid = 21'b000011010111100001101;
		14'b11101000111001:	sigmoid = 21'b000011010111111011010;
		14'b11101000111010:	sigmoid = 21'b000011011000010100111;
		14'b11101000111011:	sigmoid = 21'b000011011000101110100;
		14'b11101000111100:	sigmoid = 21'b000011011001001000001;
		14'b11101000111101:	sigmoid = 21'b000011011001100001111;
		14'b11101000111110:	sigmoid = 21'b000011011001111011101;
		14'b11101000111111:	sigmoid = 21'b000011011010010101100;
		14'b11101001000000:	sigmoid = 21'b000011011010101111010;
		14'b11101001000001:	sigmoid = 21'b000011011011001001010;
		14'b11101001000010:	sigmoid = 21'b000011011011100011001;
		14'b11101001000011:	sigmoid = 21'b000011011011111101001;
		14'b11101001000100:	sigmoid = 21'b000011011100010111010;
		14'b11101001000101:	sigmoid = 21'b000011011100110001010;
		14'b11101001000110:	sigmoid = 21'b000011011101001011011;
		14'b11101001000111:	sigmoid = 21'b000011011101100101101;
		14'b11101001001000:	sigmoid = 21'b000011011101111111110;
		14'b11101001001001:	sigmoid = 21'b000011011110011010001;
		14'b11101001001010:	sigmoid = 21'b000011011110110100011;
		14'b11101001001011:	sigmoid = 21'b000011011111001110110;
		14'b11101001001100:	sigmoid = 21'b000011011111101001001;
		14'b11101001001101:	sigmoid = 21'b000011100000000011101;
		14'b11101001001110:	sigmoid = 21'b000011100000011110001;
		14'b11101001001111:	sigmoid = 21'b000011100000111000101;
		14'b11101001010000:	sigmoid = 21'b000011100001010011010;
		14'b11101001010001:	sigmoid = 21'b000011100001101101111;
		14'b11101001010010:	sigmoid = 21'b000011100010001000101;
		14'b11101001010011:	sigmoid = 21'b000011100010100011010;
		14'b11101001010100:	sigmoid = 21'b000011100010111110001;
		14'b11101001010101:	sigmoid = 21'b000011100011011000111;
		14'b11101001010110:	sigmoid = 21'b000011100011110011110;
		14'b11101001010111:	sigmoid = 21'b000011100100001110101;
		14'b11101001011000:	sigmoid = 21'b000011100100101001101;
		14'b11101001011001:	sigmoid = 21'b000011100101000100101;
		14'b11101001011010:	sigmoid = 21'b000011100101011111110;
		14'b11101001011011:	sigmoid = 21'b000011100101111010110;
		14'b11101001011100:	sigmoid = 21'b000011100110010110000;
		14'b11101001011101:	sigmoid = 21'b000011100110110001001;
		14'b11101001011110:	sigmoid = 21'b000011100111001100011;
		14'b11101001011111:	sigmoid = 21'b000011100111100111110;
		14'b11101001100000:	sigmoid = 21'b000011101000000011000;
		14'b11101001100001:	sigmoid = 21'b000011101000011110011;
		14'b11101001100010:	sigmoid = 21'b000011101000111001111;
		14'b11101001100011:	sigmoid = 21'b000011101001010101011;
		14'b11101001100100:	sigmoid = 21'b000011101001110000111;
		14'b11101001100101:	sigmoid = 21'b000011101010001100100;
		14'b11101001100110:	sigmoid = 21'b000011101010101000001;
		14'b11101001100111:	sigmoid = 21'b000011101011000011110;
		14'b11101001101000:	sigmoid = 21'b000011101011011111100;
		14'b11101001101001:	sigmoid = 21'b000011101011111011010;
		14'b11101001101010:	sigmoid = 21'b000011101100010111000;
		14'b11101001101011:	sigmoid = 21'b000011101100110010111;
		14'b11101001101100:	sigmoid = 21'b000011101101001110111;
		14'b11101001101101:	sigmoid = 21'b000011101101101010110;
		14'b11101001101110:	sigmoid = 21'b000011101110000110110;
		14'b11101001101111:	sigmoid = 21'b000011101110100010111;
		14'b11101001110000:	sigmoid = 21'b000011101110111111000;
		14'b11101001110001:	sigmoid = 21'b000011101111011011001;
		14'b11101001110010:	sigmoid = 21'b000011101111110111010;
		14'b11101001110011:	sigmoid = 21'b000011110000010011100;
		14'b11101001110100:	sigmoid = 21'b000011110000101111111;
		14'b11101001110101:	sigmoid = 21'b000011110001001100010;
		14'b11101001110110:	sigmoid = 21'b000011110001101000101;
		14'b11101001110111:	sigmoid = 21'b000011110010000101000;
		14'b11101001111000:	sigmoid = 21'b000011110010100001100;
		14'b11101001111001:	sigmoid = 21'b000011110010111110001;
		14'b11101001111010:	sigmoid = 21'b000011110011011010110;
		14'b11101001111011:	sigmoid = 21'b000011110011110111011;
		14'b11101001111100:	sigmoid = 21'b000011110100010100000;
		14'b11101001111101:	sigmoid = 21'b000011110100110000110;
		14'b11101001111110:	sigmoid = 21'b000011110101001101100;
		14'b11101001111111:	sigmoid = 21'b000011110101101010011;
		14'b11101010000000:	sigmoid = 21'b000011110110000111010;
		14'b11101010000001:	sigmoid = 21'b000011110110100100010;
		14'b11101010000010:	sigmoid = 21'b000011110111000001010;
		14'b11101010000011:	sigmoid = 21'b000011110111011110010;
		14'b11101010000100:	sigmoid = 21'b000011110111111011011;
		14'b11101010000101:	sigmoid = 21'b000011111000011000100;
		14'b11101010000110:	sigmoid = 21'b000011111000110101101;
		14'b11101010000111:	sigmoid = 21'b000011111001010010111;
		14'b11101010001000:	sigmoid = 21'b000011111001110000010;
		14'b11101010001001:	sigmoid = 21'b000011111010001101100;
		14'b11101010001010:	sigmoid = 21'b000011111010101011000;
		14'b11101010001011:	sigmoid = 21'b000011111011001000011;
		14'b11101010001100:	sigmoid = 21'b000011111011100101111;
		14'b11101010001101:	sigmoid = 21'b000011111100000011011;
		14'b11101010001110:	sigmoid = 21'b000011111100100001000;
		14'b11101010001111:	sigmoid = 21'b000011111100111110101;
		14'b11101010010000:	sigmoid = 21'b000011111101011100011;
		14'b11101010010001:	sigmoid = 21'b000011111101111010001;
		14'b11101010010010:	sigmoid = 21'b000011111110010111111;
		14'b11101010010011:	sigmoid = 21'b000011111110110101110;
		14'b11101010010100:	sigmoid = 21'b000011111111010011101;
		14'b11101010010101:	sigmoid = 21'b000011111111110001101;
		14'b11101010010110:	sigmoid = 21'b000100000000001111101;
		14'b11101010010111:	sigmoid = 21'b000100000000101101101;
		14'b11101010011000:	sigmoid = 21'b000100000001001011110;
		14'b11101010011001:	sigmoid = 21'b000100000001101001111;
		14'b11101010011010:	sigmoid = 21'b000100000010001000001;
		14'b11101010011011:	sigmoid = 21'b000100000010100110011;
		14'b11101010011100:	sigmoid = 21'b000100000011000100101;
		14'b11101010011101:	sigmoid = 21'b000100000011100011000;
		14'b11101010011110:	sigmoid = 21'b000100000100000001100;
		14'b11101010011111:	sigmoid = 21'b000100000100011111111;
		14'b11101010100000:	sigmoid = 21'b000100000100111110100;
		14'b11101010100001:	sigmoid = 21'b000100000101011101000;
		14'b11101010100010:	sigmoid = 21'b000100000101111011101;
		14'b11101010100011:	sigmoid = 21'b000100000110011010010;
		14'b11101010100100:	sigmoid = 21'b000100000110111001000;
		14'b11101010100101:	sigmoid = 21'b000100000111010111110;
		14'b11101010100110:	sigmoid = 21'b000100000111110110101;
		14'b11101010100111:	sigmoid = 21'b000100001000010101100;
		14'b11101010101000:	sigmoid = 21'b000100001000110100100;
		14'b11101010101001:	sigmoid = 21'b000100001001010011100;
		14'b11101010101010:	sigmoid = 21'b000100001001110010100;
		14'b11101010101011:	sigmoid = 21'b000100001010010001101;
		14'b11101010101100:	sigmoid = 21'b000100001010110000110;
		14'b11101010101101:	sigmoid = 21'b000100001011001111111;
		14'b11101010101110:	sigmoid = 21'b000100001011101111001;
		14'b11101010101111:	sigmoid = 21'b000100001100001110100;
		14'b11101010110000:	sigmoid = 21'b000100001100101101111;
		14'b11101010110001:	sigmoid = 21'b000100001101001101010;
		14'b11101010110010:	sigmoid = 21'b000100001101101100110;
		14'b11101010110011:	sigmoid = 21'b000100001110001100010;
		14'b11101010110100:	sigmoid = 21'b000100001110101011111;
		14'b11101010110101:	sigmoid = 21'b000100001111001011100;
		14'b11101010110110:	sigmoid = 21'b000100001111101011001;
		14'b11101010110111:	sigmoid = 21'b000100010000001010111;
		14'b11101010111000:	sigmoid = 21'b000100010000101010101;
		14'b11101010111001:	sigmoid = 21'b000100010001001010100;
		14'b11101010111010:	sigmoid = 21'b000100010001101010011;
		14'b11101010111011:	sigmoid = 21'b000100010010001010011;
		14'b11101010111100:	sigmoid = 21'b000100010010101010011;
		14'b11101010111101:	sigmoid = 21'b000100010011001010011;
		14'b11101010111110:	sigmoid = 21'b000100010011101010100;
		14'b11101010111111:	sigmoid = 21'b000100010100001010101;
		14'b11101011000000:	sigmoid = 21'b000100010100101010111;
		14'b11101011000001:	sigmoid = 21'b000100010101001011001;
		14'b11101011000010:	sigmoid = 21'b000100010101101011100;
		14'b11101011000011:	sigmoid = 21'b000100010110001011111;
		14'b11101011000100:	sigmoid = 21'b000100010110101100011;
		14'b11101011000101:	sigmoid = 21'b000100010111001100111;
		14'b11101011000110:	sigmoid = 21'b000100010111101101011;
		14'b11101011000111:	sigmoid = 21'b000100011000001110000;
		14'b11101011001000:	sigmoid = 21'b000100011000101110101;
		14'b11101011001001:	sigmoid = 21'b000100011001001111011;
		14'b11101011001010:	sigmoid = 21'b000100011001110000001;
		14'b11101011001011:	sigmoid = 21'b000100011010010000111;
		14'b11101011001100:	sigmoid = 21'b000100011010110001111;
		14'b11101011001101:	sigmoid = 21'b000100011011010010110;
		14'b11101011001110:	sigmoid = 21'b000100011011110011110;
		14'b11101011001111:	sigmoid = 21'b000100011100010100110;
		14'b11101011010000:	sigmoid = 21'b000100011100110101111;
		14'b11101011010001:	sigmoid = 21'b000100011101010111000;
		14'b11101011010010:	sigmoid = 21'b000100011101111000010;
		14'b11101011010011:	sigmoid = 21'b000100011110011001100;
		14'b11101011010100:	sigmoid = 21'b000100011110111010111;
		14'b11101011010101:	sigmoid = 21'b000100011111011100010;
		14'b11101011010110:	sigmoid = 21'b000100011111111101101;
		14'b11101011010111:	sigmoid = 21'b000100100000011111001;
		14'b11101011011000:	sigmoid = 21'b000100100001000000110;
		14'b11101011011001:	sigmoid = 21'b000100100001100010011;
		14'b11101011011010:	sigmoid = 21'b000100100010000100000;
		14'b11101011011011:	sigmoid = 21'b000100100010100101110;
		14'b11101011011100:	sigmoid = 21'b000100100011000111100;
		14'b11101011011101:	sigmoid = 21'b000100100011101001010;
		14'b11101011011110:	sigmoid = 21'b000100100100001011010;
		14'b11101011011111:	sigmoid = 21'b000100100100101101001;
		14'b11101011100000:	sigmoid = 21'b000100100101001111001;
		14'b11101011100001:	sigmoid = 21'b000100100101110001010;
		14'b11101011100010:	sigmoid = 21'b000100100110010011011;
		14'b11101011100011:	sigmoid = 21'b000100100110110101100;
		14'b11101011100100:	sigmoid = 21'b000100100111010111110;
		14'b11101011100101:	sigmoid = 21'b000100100111111010000;
		14'b11101011100110:	sigmoid = 21'b000100101000011100011;
		14'b11101011100111:	sigmoid = 21'b000100101000111110110;
		14'b11101011101000:	sigmoid = 21'b000100101001100001010;
		14'b11101011101001:	sigmoid = 21'b000100101010000011110;
		14'b11101011101010:	sigmoid = 21'b000100101010100110010;
		14'b11101011101011:	sigmoid = 21'b000100101011001001000;
		14'b11101011101100:	sigmoid = 21'b000100101011101011101;
		14'b11101011101101:	sigmoid = 21'b000100101100001110011;
		14'b11101011101110:	sigmoid = 21'b000100101100110001001;
		14'b11101011101111:	sigmoid = 21'b000100101101010100000;
		14'b11101011110000:	sigmoid = 21'b000100101101110111000;
		14'b11101011110001:	sigmoid = 21'b000100101110011010000;
		14'b11101011110010:	sigmoid = 21'b000100101110111101000;
		14'b11101011110011:	sigmoid = 21'b000100101111100000001;
		14'b11101011110100:	sigmoid = 21'b000100110000000011010;
		14'b11101011110101:	sigmoid = 21'b000100110000100110100;
		14'b11101011110110:	sigmoid = 21'b000100110001001001110;
		14'b11101011110111:	sigmoid = 21'b000100110001101101001;
		14'b11101011111000:	sigmoid = 21'b000100110010010000100;
		14'b11101011111001:	sigmoid = 21'b000100110010110011111;
		14'b11101011111010:	sigmoid = 21'b000100110011010111011;
		14'b11101011111011:	sigmoid = 21'b000100110011111011000;
		14'b11101011111100:	sigmoid = 21'b000100110100011110101;
		14'b11101011111101:	sigmoid = 21'b000100110101000010010;
		14'b11101011111110:	sigmoid = 21'b000100110101100110000;
		14'b11101011111111:	sigmoid = 21'b000100110110001001111;
		14'b11101100000000:	sigmoid = 21'b000100110110101101110;
		14'b11101100000001:	sigmoid = 21'b000100110111010001101;
		14'b11101100000010:	sigmoid = 21'b000100110111110101101;
		14'b11101100000011:	sigmoid = 21'b000100111000011001101;
		14'b11101100000100:	sigmoid = 21'b000100111000111101110;
		14'b11101100000101:	sigmoid = 21'b000100111001100001111;
		14'b11101100000110:	sigmoid = 21'b000100111010000110001;
		14'b11101100000111:	sigmoid = 21'b000100111010101010011;
		14'b11101100001000:	sigmoid = 21'b000100111011001110110;
		14'b11101100001001:	sigmoid = 21'b000100111011110011001;
		14'b11101100001010:	sigmoid = 21'b000100111100010111101;
		14'b11101100001011:	sigmoid = 21'b000100111100111100001;
		14'b11101100001100:	sigmoid = 21'b000100111101100000110;
		14'b11101100001101:	sigmoid = 21'b000100111110000101011;
		14'b11101100001110:	sigmoid = 21'b000100111110101010001;
		14'b11101100001111:	sigmoid = 21'b000100111111001110111;
		14'b11101100010000:	sigmoid = 21'b000100111111110011101;
		14'b11101100010001:	sigmoid = 21'b000101000000011000100;
		14'b11101100010010:	sigmoid = 21'b000101000000111101100;
		14'b11101100010011:	sigmoid = 21'b000101000001100010100;
		14'b11101100010100:	sigmoid = 21'b000101000010000111101;
		14'b11101100010101:	sigmoid = 21'b000101000010101100110;
		14'b11101100010110:	sigmoid = 21'b000101000011010001111;
		14'b11101100010111:	sigmoid = 21'b000101000011110111001;
		14'b11101100011000:	sigmoid = 21'b000101000100011100100;
		14'b11101100011001:	sigmoid = 21'b000101000101000001111;
		14'b11101100011010:	sigmoid = 21'b000101000101100111010;
		14'b11101100011011:	sigmoid = 21'b000101000110001100110;
		14'b11101100011100:	sigmoid = 21'b000101000110110010011;
		14'b11101100011101:	sigmoid = 21'b000101000111010111111;
		14'b11101100011110:	sigmoid = 21'b000101000111111101101;
		14'b11101100011111:	sigmoid = 21'b000101001000100011011;
		14'b11101100100000:	sigmoid = 21'b000101001001001001001;
		14'b11101100100001:	sigmoid = 21'b000101001001101111000;
		14'b11101100100010:	sigmoid = 21'b000101001010010101000;
		14'b11101100100011:	sigmoid = 21'b000101001010111011000;
		14'b11101100100100:	sigmoid = 21'b000101001011100001000;
		14'b11101100100101:	sigmoid = 21'b000101001100000111001;
		14'b11101100100110:	sigmoid = 21'b000101001100101101010;
		14'b11101100100111:	sigmoid = 21'b000101001101010011100;
		14'b11101100101000:	sigmoid = 21'b000101001101111001111;
		14'b11101100101001:	sigmoid = 21'b000101001110100000010;
		14'b11101100101010:	sigmoid = 21'b000101001111000110101;
		14'b11101100101011:	sigmoid = 21'b000101001111101101001;
		14'b11101100101100:	sigmoid = 21'b000101010000010011110;
		14'b11101100101101:	sigmoid = 21'b000101010000111010011;
		14'b11101100101110:	sigmoid = 21'b000101010001100001000;
		14'b11101100101111:	sigmoid = 21'b000101010010000111110;
		14'b11101100110000:	sigmoid = 21'b000101010010101110100;
		14'b11101100110001:	sigmoid = 21'b000101010011010101011;
		14'b11101100110010:	sigmoid = 21'b000101010011111100011;
		14'b11101100110011:	sigmoid = 21'b000101010100100011011;
		14'b11101100110100:	sigmoid = 21'b000101010101001010011;
		14'b11101100110101:	sigmoid = 21'b000101010101110001100;
		14'b11101100110110:	sigmoid = 21'b000101010110011000110;
		14'b11101100110111:	sigmoid = 21'b000101010111000000000;
		14'b11101100111000:	sigmoid = 21'b000101010111100111010;
		14'b11101100111001:	sigmoid = 21'b000101011000001110101;
		14'b11101100111010:	sigmoid = 21'b000101011000110110001;
		14'b11101100111011:	sigmoid = 21'b000101011001011101101;
		14'b11101100111100:	sigmoid = 21'b000101011010000101010;
		14'b11101100111101:	sigmoid = 21'b000101011010101100111;
		14'b11101100111110:	sigmoid = 21'b000101011011010100100;
		14'b11101100111111:	sigmoid = 21'b000101011011111100010;
		14'b11101101000000:	sigmoid = 21'b000101011100100100001;
		14'b11101101000001:	sigmoid = 21'b000101011101001100000;
		14'b11101101000010:	sigmoid = 21'b000101011101110100000;
		14'b11101101000011:	sigmoid = 21'b000101011110011100000;
		14'b11101101000100:	sigmoid = 21'b000101011111000100001;
		14'b11101101000101:	sigmoid = 21'b000101011111101100010;
		14'b11101101000110:	sigmoid = 21'b000101100000010100100;
		14'b11101101000111:	sigmoid = 21'b000101100000111100110;
		14'b11101101001000:	sigmoid = 21'b000101100001100101001;
		14'b11101101001001:	sigmoid = 21'b000101100010001101100;
		14'b11101101001010:	sigmoid = 21'b000101100010110110000;
		14'b11101101001011:	sigmoid = 21'b000101100011011110100;
		14'b11101101001100:	sigmoid = 21'b000101100100000111001;
		14'b11101101001101:	sigmoid = 21'b000101100100101111111;
		14'b11101101001110:	sigmoid = 21'b000101100101011000101;
		14'b11101101001111:	sigmoid = 21'b000101100110000001011;
		14'b11101101010000:	sigmoid = 21'b000101100110101010010;
		14'b11101101010001:	sigmoid = 21'b000101100111010011010;
		14'b11101101010010:	sigmoid = 21'b000101100111111100010;
		14'b11101101010011:	sigmoid = 21'b000101101000100101010;
		14'b11101101010100:	sigmoid = 21'b000101101001001110011;
		14'b11101101010101:	sigmoid = 21'b000101101001110111101;
		14'b11101101010110:	sigmoid = 21'b000101101010100000111;
		14'b11101101010111:	sigmoid = 21'b000101101011001010010;
		14'b11101101011000:	sigmoid = 21'b000101101011110011101;
		14'b11101101011001:	sigmoid = 21'b000101101100011101001;
		14'b11101101011010:	sigmoid = 21'b000101101101000110101;
		14'b11101101011011:	sigmoid = 21'b000101101101110000010;
		14'b11101101011100:	sigmoid = 21'b000101101110011001111;
		14'b11101101011101:	sigmoid = 21'b000101101111000011101;
		14'b11101101011110:	sigmoid = 21'b000101101111101101100;
		14'b11101101011111:	sigmoid = 21'b000101110000010111011;
		14'b11101101100000:	sigmoid = 21'b000101110001000001010;
		14'b11101101100001:	sigmoid = 21'b000101110001101011010;
		14'b11101101100010:	sigmoid = 21'b000101110010010101011;
		14'b11101101100011:	sigmoid = 21'b000101110010111111100;
		14'b11101101100100:	sigmoid = 21'b000101110011101001110;
		14'b11101101100101:	sigmoid = 21'b000101110100010100000;
		14'b11101101100110:	sigmoid = 21'b000101110100111110011;
		14'b11101101100111:	sigmoid = 21'b000101110101101000110;
		14'b11101101101000:	sigmoid = 21'b000101110110010011010;
		14'b11101101101001:	sigmoid = 21'b000101110110111101110;
		14'b11101101101010:	sigmoid = 21'b000101110111101000011;
		14'b11101101101011:	sigmoid = 21'b000101111000010011000;
		14'b11101101101100:	sigmoid = 21'b000101111000111101110;
		14'b11101101101101:	sigmoid = 21'b000101111001101000101;
		14'b11101101101110:	sigmoid = 21'b000101111010010011100;
		14'b11101101101111:	sigmoid = 21'b000101111010111110100;
		14'b11101101110000:	sigmoid = 21'b000101111011101001100;
		14'b11101101110001:	sigmoid = 21'b000101111100010100101;
		14'b11101101110010:	sigmoid = 21'b000101111100111111110;
		14'b11101101110011:	sigmoid = 21'b000101111101101011000;
		14'b11101101110100:	sigmoid = 21'b000101111110010110010;
		14'b11101101110101:	sigmoid = 21'b000101111111000001101;
		14'b11101101110110:	sigmoid = 21'b000101111111101101001;
		14'b11101101110111:	sigmoid = 21'b000110000000011000101;
		14'b11101101111000:	sigmoid = 21'b000110000001000100001;
		14'b11101101111001:	sigmoid = 21'b000110000001101111110;
		14'b11101101111010:	sigmoid = 21'b000110000010011011100;
		14'b11101101111011:	sigmoid = 21'b000110000011000111010;
		14'b11101101111100:	sigmoid = 21'b000110000011110011001;
		14'b11101101111101:	sigmoid = 21'b000110000100011111000;
		14'b11101101111110:	sigmoid = 21'b000110000101001011000;
		14'b11101101111111:	sigmoid = 21'b000110000101110111001;
		14'b11101110000000:	sigmoid = 21'b000110000110100011010;
		14'b11101110000001:	sigmoid = 21'b000110000111001111011;
		14'b11101110000010:	sigmoid = 21'b000110000111111011110;
		14'b11101110000011:	sigmoid = 21'b000110001000101000000;
		14'b11101110000100:	sigmoid = 21'b000110001001010100100;
		14'b11101110000101:	sigmoid = 21'b000110001010000000111;
		14'b11101110000110:	sigmoid = 21'b000110001010101101100;
		14'b11101110000111:	sigmoid = 21'b000110001011011010001;
		14'b11101110001000:	sigmoid = 21'b000110001100000110110;
		14'b11101110001001:	sigmoid = 21'b000110001100110011100;
		14'b11101110001010:	sigmoid = 21'b000110001101100000011;
		14'b11101110001011:	sigmoid = 21'b000110001110001101010;
		14'b11101110001100:	sigmoid = 21'b000110001110111010010;
		14'b11101110001101:	sigmoid = 21'b000110001111100111010;
		14'b11101110001110:	sigmoid = 21'b000110010000010100011;
		14'b11101110001111:	sigmoid = 21'b000110010001000001101;
		14'b11101110010000:	sigmoid = 21'b000110010001101110111;
		14'b11101110010001:	sigmoid = 21'b000110010010011100001;
		14'b11101110010010:	sigmoid = 21'b000110010011001001101;
		14'b11101110010011:	sigmoid = 21'b000110010011110111000;
		14'b11101110010100:	sigmoid = 21'b000110010100100100101;
		14'b11101110010101:	sigmoid = 21'b000110010101010010010;
		14'b11101110010110:	sigmoid = 21'b000110010101111111111;
		14'b11101110010111:	sigmoid = 21'b000110010110101101101;
		14'b11101110011000:	sigmoid = 21'b000110010111011011100;
		14'b11101110011001:	sigmoid = 21'b000110011000001001011;
		14'b11101110011010:	sigmoid = 21'b000110011000110111011;
		14'b11101110011011:	sigmoid = 21'b000110011001100101011;
		14'b11101110011100:	sigmoid = 21'b000110011010010011100;
		14'b11101110011101:	sigmoid = 21'b000110011011000001101;
		14'b11101110011110:	sigmoid = 21'b000110011011101111111;
		14'b11101110011111:	sigmoid = 21'b000110011100011110010;
		14'b11101110100000:	sigmoid = 21'b000110011101001100101;
		14'b11101110100001:	sigmoid = 21'b000110011101111011001;
		14'b11101110100010:	sigmoid = 21'b000110011110101001101;
		14'b11101110100011:	sigmoid = 21'b000110011111011000010;
		14'b11101110100100:	sigmoid = 21'b000110100000000111000;
		14'b11101110100101:	sigmoid = 21'b000110100000110101110;
		14'b11101110100110:	sigmoid = 21'b000110100001100100101;
		14'b11101110100111:	sigmoid = 21'b000110100010010011100;
		14'b11101110101000:	sigmoid = 21'b000110100011000010100;
		14'b11101110101001:	sigmoid = 21'b000110100011110001100;
		14'b11101110101010:	sigmoid = 21'b000110100100100000110;
		14'b11101110101011:	sigmoid = 21'b000110100101001111111;
		14'b11101110101100:	sigmoid = 21'b000110100101111111001;
		14'b11101110101101:	sigmoid = 21'b000110100110101110100;
		14'b11101110101110:	sigmoid = 21'b000110100111011110000;
		14'b11101110101111:	sigmoid = 21'b000110101000001101100;
		14'b11101110110000:	sigmoid = 21'b000110101000111101000;
		14'b11101110110001:	sigmoid = 21'b000110101001101100101;
		14'b11101110110010:	sigmoid = 21'b000110101010011100011;
		14'b11101110110011:	sigmoid = 21'b000110101011001100001;
		14'b11101110110100:	sigmoid = 21'b000110101011111100000;
		14'b11101110110101:	sigmoid = 21'b000110101100101100000;
		14'b11101110110110:	sigmoid = 21'b000110101101011100000;
		14'b11101110110111:	sigmoid = 21'b000110101110001100001;
		14'b11101110111000:	sigmoid = 21'b000110101110111100010;
		14'b11101110111001:	sigmoid = 21'b000110101111101100100;
		14'b11101110111010:	sigmoid = 21'b000110110000011100110;
		14'b11101110111011:	sigmoid = 21'b000110110001001101001;
		14'b11101110111100:	sigmoid = 21'b000110110001111101101;
		14'b11101110111101:	sigmoid = 21'b000110110010101110001;
		14'b11101110111110:	sigmoid = 21'b000110110011011110110;
		14'b11101110111111:	sigmoid = 21'b000110110100001111100;
		14'b11101111000000:	sigmoid = 21'b000110110101000000010;
		14'b11101111000001:	sigmoid = 21'b000110110101110001001;
		14'b11101111000010:	sigmoid = 21'b000110110110100010000;
		14'b11101111000011:	sigmoid = 21'b000110110111010011000;
		14'b11101111000100:	sigmoid = 21'b000110111000000100000;
		14'b11101111000101:	sigmoid = 21'b000110111000110101001;
		14'b11101111000110:	sigmoid = 21'b000110111001100110011;
		14'b11101111000111:	sigmoid = 21'b000110111010010111101;
		14'b11101111001000:	sigmoid = 21'b000110111011001001000;
		14'b11101111001001:	sigmoid = 21'b000110111011111010100;
		14'b11101111001010:	sigmoid = 21'b000110111100101100000;
		14'b11101111001011:	sigmoid = 21'b000110111101011101101;
		14'b11101111001100:	sigmoid = 21'b000110111110001111010;
		14'b11101111001101:	sigmoid = 21'b000110111111000001000;
		14'b11101111001110:	sigmoid = 21'b000110111111110010110;
		14'b11101111001111:	sigmoid = 21'b000111000000100100101;
		14'b11101111010000:	sigmoid = 21'b000111000001010110101;
		14'b11101111010001:	sigmoid = 21'b000111000010001000110;
		14'b11101111010010:	sigmoid = 21'b000111000010111010111;
		14'b11101111010011:	sigmoid = 21'b000111000011101101000;
		14'b11101111010100:	sigmoid = 21'b000111000100011111010;
		14'b11101111010101:	sigmoid = 21'b000111000101010001101;
		14'b11101111010110:	sigmoid = 21'b000111000110000100001;
		14'b11101111010111:	sigmoid = 21'b000111000110110110101;
		14'b11101111011000:	sigmoid = 21'b000111000111101001001;
		14'b11101111011001:	sigmoid = 21'b000111001000011011110;
		14'b11101111011010:	sigmoid = 21'b000111001001001110100;
		14'b11101111011011:	sigmoid = 21'b000111001010000001011;
		14'b11101111011100:	sigmoid = 21'b000111001010110100010;
		14'b11101111011101:	sigmoid = 21'b000111001011100111010;
		14'b11101111011110:	sigmoid = 21'b000111001100011010010;
		14'b11101111011111:	sigmoid = 21'b000111001101001101011;
		14'b11101111100000:	sigmoid = 21'b000111001110000000101;
		14'b11101111100001:	sigmoid = 21'b000111001110110011111;
		14'b11101111100010:	sigmoid = 21'b000111001111100111010;
		14'b11101111100011:	sigmoid = 21'b000111010000011010101;
		14'b11101111100100:	sigmoid = 21'b000111010001001110001;
		14'b11101111100101:	sigmoid = 21'b000111010010000001110;
		14'b11101111100110:	sigmoid = 21'b000111010010110101011;
		14'b11101111100111:	sigmoid = 21'b000111010011101001001;
		14'b11101111101000:	sigmoid = 21'b000111010100011101000;
		14'b11101111101001:	sigmoid = 21'b000111010101010000111;
		14'b11101111101010:	sigmoid = 21'b000111010110000100111;
		14'b11101111101011:	sigmoid = 21'b000111010110111000111;
		14'b11101111101100:	sigmoid = 21'b000111010111101101000;
		14'b11101111101101:	sigmoid = 21'b000111011000100001010;
		14'b11101111101110:	sigmoid = 21'b000111011001010101100;
		14'b11101111101111:	sigmoid = 21'b000111011010001001111;
		14'b11101111110000:	sigmoid = 21'b000111011010111110011;
		14'b11101111110001:	sigmoid = 21'b000111011011110010111;
		14'b11101111110010:	sigmoid = 21'b000111011100100111100;
		14'b11101111110011:	sigmoid = 21'b000111011101011100001;
		14'b11101111110100:	sigmoid = 21'b000111011110010000111;
		14'b11101111110101:	sigmoid = 21'b000111011111000101110;
		14'b11101111110110:	sigmoid = 21'b000111011111111010101;
		14'b11101111110111:	sigmoid = 21'b000111100000101111101;
		14'b11101111111000:	sigmoid = 21'b000111100001100100110;
		14'b11101111111001:	sigmoid = 21'b000111100010011001111;
		14'b11101111111010:	sigmoid = 21'b000111100011001111001;
		14'b11101111111011:	sigmoid = 21'b000111100100000100100;
		14'b11101111111100:	sigmoid = 21'b000111100100111001111;
		14'b11101111111101:	sigmoid = 21'b000111100101101111011;
		14'b11101111111110:	sigmoid = 21'b000111100110100100111;
		14'b11101111111111:	sigmoid = 21'b000111100111011010100;
		14'b11110000000000:	sigmoid = 21'b000111101000010000010;
		14'b11110000000001:	sigmoid = 21'b000111101001000110001;
		14'b11110000000010:	sigmoid = 21'b000111101001111100000;
		14'b11110000000011:	sigmoid = 21'b000111101010110001111;
		14'b11110000000100:	sigmoid = 21'b000111101011100111111;
		14'b11110000000101:	sigmoid = 21'b000111101100011110000;
		14'b11110000000110:	sigmoid = 21'b000111101101010100010;
		14'b11110000000111:	sigmoid = 21'b000111101110001010100;
		14'b11110000001000:	sigmoid = 21'b000111101111000000111;
		14'b11110000001001:	sigmoid = 21'b000111101111110111011;
		14'b11110000001010:	sigmoid = 21'b000111110000101101111;
		14'b11110000001011:	sigmoid = 21'b000111110001100100100;
		14'b11110000001100:	sigmoid = 21'b000111110010011011001;
		14'b11110000001101:	sigmoid = 21'b000111110011010001111;
		14'b11110000001110:	sigmoid = 21'b000111110100001000110;
		14'b11110000001111:	sigmoid = 21'b000111110100111111101;
		14'b11110000010000:	sigmoid = 21'b000111110101110110101;
		14'b11110000010001:	sigmoid = 21'b000111110110101101110;
		14'b11110000010010:	sigmoid = 21'b000111110111100100111;
		14'b11110000010011:	sigmoid = 21'b000111111000011100001;
		14'b11110000010100:	sigmoid = 21'b000111111001010011100;
		14'b11110000010101:	sigmoid = 21'b000111111010001010111;
		14'b11110000010110:	sigmoid = 21'b000111111011000010011;
		14'b11110000010111:	sigmoid = 21'b000111111011111010000;
		14'b11110000011000:	sigmoid = 21'b000111111100110001101;
		14'b11110000011001:	sigmoid = 21'b000111111101101001011;
		14'b11110000011010:	sigmoid = 21'b000111111110100001010;
		14'b11110000011011:	sigmoid = 21'b000111111111011001001;
		14'b11110000011100:	sigmoid = 21'b001000000000010001001;
		14'b11110000011101:	sigmoid = 21'b001000000001001001001;
		14'b11110000011110:	sigmoid = 21'b001000000010000001010;
		14'b11110000011111:	sigmoid = 21'b001000000010111001100;
		14'b11110000100000:	sigmoid = 21'b001000000011110001111;
		14'b11110000100001:	sigmoid = 21'b001000000100101010010;
		14'b11110000100010:	sigmoid = 21'b001000000101100010110;
		14'b11110000100011:	sigmoid = 21'b001000000110011011010;
		14'b11110000100100:	sigmoid = 21'b001000000111010011111;
		14'b11110000100101:	sigmoid = 21'b001000001000001100101;
		14'b11110000100110:	sigmoid = 21'b001000001001000101100;
		14'b11110000100111:	sigmoid = 21'b001000001001111110011;
		14'b11110000101000:	sigmoid = 21'b001000001010110111010;
		14'b11110000101001:	sigmoid = 21'b001000001011110000011;
		14'b11110000101010:	sigmoid = 21'b001000001100101001100;
		14'b11110000101011:	sigmoid = 21'b001000001101100010110;
		14'b11110000101100:	sigmoid = 21'b001000001110011100000;
		14'b11110000101101:	sigmoid = 21'b001000001111010101011;
		14'b11110000101110:	sigmoid = 21'b001000010000001110111;
		14'b11110000101111:	sigmoid = 21'b001000010001001000100;
		14'b11110000110000:	sigmoid = 21'b001000010010000010001;
		14'b11110000110001:	sigmoid = 21'b001000010010111011110;
		14'b11110000110010:	sigmoid = 21'b001000010011110101101;
		14'b11110000110011:	sigmoid = 21'b001000010100101111100;
		14'b11110000110100:	sigmoid = 21'b001000010101101001100;
		14'b11110000110101:	sigmoid = 21'b001000010110100011100;
		14'b11110000110110:	sigmoid = 21'b001000010111011101101;
		14'b11110000110111:	sigmoid = 21'b001000011000010111111;
		14'b11110000111000:	sigmoid = 21'b001000011001010010010;
		14'b11110000111001:	sigmoid = 21'b001000011010001100101;
		14'b11110000111010:	sigmoid = 21'b001000011011000111001;
		14'b11110000111011:	sigmoid = 21'b001000011100000001101;
		14'b11110000111100:	sigmoid = 21'b001000011100111100010;
		14'b11110000111101:	sigmoid = 21'b001000011101110111000;
		14'b11110000111110:	sigmoid = 21'b001000011110110001111;
		14'b11110000111111:	sigmoid = 21'b001000011111101100110;
		14'b11110001000000:	sigmoid = 21'b001000100000100111110;
		14'b11110001000001:	sigmoid = 21'b001000100001100010110;
		14'b11110001000010:	sigmoid = 21'b001000100010011101111;
		14'b11110001000011:	sigmoid = 21'b001000100011011001001;
		14'b11110001000100:	sigmoid = 21'b001000100100010100100;
		14'b11110001000101:	sigmoid = 21'b001000100101001111111;
		14'b11110001000110:	sigmoid = 21'b001000100110001011011;
		14'b11110001000111:	sigmoid = 21'b001000100111000111000;
		14'b11110001001000:	sigmoid = 21'b001000101000000010101;
		14'b11110001001001:	sigmoid = 21'b001000101000111110011;
		14'b11110001001010:	sigmoid = 21'b001000101001111010010;
		14'b11110001001011:	sigmoid = 21'b001000101010110110001;
		14'b11110001001100:	sigmoid = 21'b001000101011110010001;
		14'b11110001001101:	sigmoid = 21'b001000101100101110010;
		14'b11110001001110:	sigmoid = 21'b001000101101101010011;
		14'b11110001001111:	sigmoid = 21'b001000101110100110101;
		14'b11110001010000:	sigmoid = 21'b001000101111100011000;
		14'b11110001010001:	sigmoid = 21'b001000110000011111100;
		14'b11110001010010:	sigmoid = 21'b001000110001011100000;
		14'b11110001010011:	sigmoid = 21'b001000110010011000100;
		14'b11110001010100:	sigmoid = 21'b001000110011010101010;
		14'b11110001010101:	sigmoid = 21'b001000110100010010000;
		14'b11110001010110:	sigmoid = 21'b001000110101001110111;
		14'b11110001010111:	sigmoid = 21'b001000110110001011111;
		14'b11110001011000:	sigmoid = 21'b001000110111001000111;
		14'b11110001011001:	sigmoid = 21'b001000111000000110000;
		14'b11110001011010:	sigmoid = 21'b001000111001000011010;
		14'b11110001011011:	sigmoid = 21'b001000111010000000100;
		14'b11110001011100:	sigmoid = 21'b001000111010111101111;
		14'b11110001011101:	sigmoid = 21'b001000111011111011011;
		14'b11110001011110:	sigmoid = 21'b001000111100111000111;
		14'b11110001011111:	sigmoid = 21'b001000111101110110100;
		14'b11110001100000:	sigmoid = 21'b001000111110110100010;
		14'b11110001100001:	sigmoid = 21'b001000111111110010000;
		14'b11110001100010:	sigmoid = 21'b001001000000110000000;
		14'b11110001100011:	sigmoid = 21'b001001000001101110000;
		14'b11110001100100:	sigmoid = 21'b001001000010101100000;
		14'b11110001100101:	sigmoid = 21'b001001000011101010001;
		14'b11110001100110:	sigmoid = 21'b001001000100101000011;
		14'b11110001100111:	sigmoid = 21'b001001000101100110110;
		14'b11110001101000:	sigmoid = 21'b001001000110100101001;
		14'b11110001101001:	sigmoid = 21'b001001000111100011101;
		14'b11110001101010:	sigmoid = 21'b001001001000100010010;
		14'b11110001101011:	sigmoid = 21'b001001001001100001000;
		14'b11110001101100:	sigmoid = 21'b001001001010011111110;
		14'b11110001101101:	sigmoid = 21'b001001001011011110101;
		14'b11110001101110:	sigmoid = 21'b001001001100011101100;
		14'b11110001101111:	sigmoid = 21'b001001001101011100101;
		14'b11110001110000:	sigmoid = 21'b001001001110011011110;
		14'b11110001110001:	sigmoid = 21'b001001001111011010111;
		14'b11110001110010:	sigmoid = 21'b001001010000011010010;
		14'b11110001110011:	sigmoid = 21'b001001010001011001101;
		14'b11110001110100:	sigmoid = 21'b001001010010011001000;
		14'b11110001110101:	sigmoid = 21'b001001010011011000101;
		14'b11110001110110:	sigmoid = 21'b001001010100011000010;
		14'b11110001110111:	sigmoid = 21'b001001010101011000000;
		14'b11110001111000:	sigmoid = 21'b001001010110010111111;
		14'b11110001111001:	sigmoid = 21'b001001010111010111110;
		14'b11110001111010:	sigmoid = 21'b001001011000010111110;
		14'b11110001111011:	sigmoid = 21'b001001011001010111111;
		14'b11110001111100:	sigmoid = 21'b001001011010011000000;
		14'b11110001111101:	sigmoid = 21'b001001011011011000010;
		14'b11110001111110:	sigmoid = 21'b001001011100011000101;
		14'b11110001111111:	sigmoid = 21'b001001011101011001001;
		14'b11110010000000:	sigmoid = 21'b001001011110011001101;
		14'b11110010000001:	sigmoid = 21'b001001011111011010010;
		14'b11110010000010:	sigmoid = 21'b001001100000011011000;
		14'b11110010000011:	sigmoid = 21'b001001100001011011110;
		14'b11110010000100:	sigmoid = 21'b001001100010011100101;
		14'b11110010000101:	sigmoid = 21'b001001100011011101101;
		14'b11110010000110:	sigmoid = 21'b001001100100011110110;
		14'b11110010000111:	sigmoid = 21'b001001100101011111111;
		14'b11110010001000:	sigmoid = 21'b001001100110100001001;
		14'b11110010001001:	sigmoid = 21'b001001100111100010011;
		14'b11110010001010:	sigmoid = 21'b001001101000100011111;
		14'b11110010001011:	sigmoid = 21'b001001101001100101011;
		14'b11110010001100:	sigmoid = 21'b001001101010100111000;
		14'b11110010001101:	sigmoid = 21'b001001101011101000101;
		14'b11110010001110:	sigmoid = 21'b001001101100101010100;
		14'b11110010001111:	sigmoid = 21'b001001101101101100011;
		14'b11110010010000:	sigmoid = 21'b001001101110101110010;
		14'b11110010010001:	sigmoid = 21'b001001101111110000011;
		14'b11110010010010:	sigmoid = 21'b001001110000110010100;
		14'b11110010010011:	sigmoid = 21'b001001110001110100110;
		14'b11110010010100:	sigmoid = 21'b001001110010110111000;
		14'b11110010010101:	sigmoid = 21'b001001110011111001011;
		14'b11110010010110:	sigmoid = 21'b001001110100111011111;
		14'b11110010010111:	sigmoid = 21'b001001110101111110100;
		14'b11110010011000:	sigmoid = 21'b001001110111000001010;
		14'b11110010011001:	sigmoid = 21'b001001111000000100000;
		14'b11110010011010:	sigmoid = 21'b001001111001000110111;
		14'b11110010011011:	sigmoid = 21'b001001111010001001110;
		14'b11110010011100:	sigmoid = 21'b001001111011001100111;
		14'b11110010011101:	sigmoid = 21'b001001111100010000000;
		14'b11110010011110:	sigmoid = 21'b001001111101010011001;
		14'b11110010011111:	sigmoid = 21'b001001111110010110100;
		14'b11110010100000:	sigmoid = 21'b001001111111011001111;
		14'b11110010100001:	sigmoid = 21'b001010000000011101011;
		14'b11110010100010:	sigmoid = 21'b001010000001100001000;
		14'b11110010100011:	sigmoid = 21'b001010000010100100101;
		14'b11110010100100:	sigmoid = 21'b001010000011101000011;
		14'b11110010100101:	sigmoid = 21'b001010000100101100010;
		14'b11110010100110:	sigmoid = 21'b001010000101110000010;
		14'b11110010100111:	sigmoid = 21'b001010000110110100010;
		14'b11110010101000:	sigmoid = 21'b001010000111111000011;
		14'b11110010101001:	sigmoid = 21'b001010001000111100101;
		14'b11110010101010:	sigmoid = 21'b001010001010000000111;
		14'b11110010101011:	sigmoid = 21'b001010001011000101011;
		14'b11110010101100:	sigmoid = 21'b001010001100001001111;
		14'b11110010101101:	sigmoid = 21'b001010001101001110011;
		14'b11110010101110:	sigmoid = 21'b001010001110010011001;
		14'b11110010101111:	sigmoid = 21'b001010001111010111111;
		14'b11110010110000:	sigmoid = 21'b001010010000011100110;
		14'b11110010110001:	sigmoid = 21'b001010010001100001101;
		14'b11110010110010:	sigmoid = 21'b001010010010100110110;
		14'b11110010110011:	sigmoid = 21'b001010010011101011111;
		14'b11110010110100:	sigmoid = 21'b001010010100110001001;
		14'b11110010110101:	sigmoid = 21'b001010010101110110011;
		14'b11110010110110:	sigmoid = 21'b001010010110111011110;
		14'b11110010110111:	sigmoid = 21'b001010011000000001010;
		14'b11110010111000:	sigmoid = 21'b001010011001000110111;
		14'b11110010111001:	sigmoid = 21'b001010011010001100101;
		14'b11110010111010:	sigmoid = 21'b001010011011010010011;
		14'b11110010111011:	sigmoid = 21'b001010011100011000010;
		14'b11110010111100:	sigmoid = 21'b001010011101011110001;
		14'b11110010111101:	sigmoid = 21'b001010011110100100010;
		14'b11110010111110:	sigmoid = 21'b001010011111101010011;
		14'b11110010111111:	sigmoid = 21'b001010100000110000101;
		14'b11110011000000:	sigmoid = 21'b001010100001110111000;
		14'b11110011000001:	sigmoid = 21'b001010100010111101011;
		14'b11110011000010:	sigmoid = 21'b001010100100000011111;
		14'b11110011000011:	sigmoid = 21'b001010100101001010100;
		14'b11110011000100:	sigmoid = 21'b001010100110010001001;
		14'b11110011000101:	sigmoid = 21'b001010100111011000000;
		14'b11110011000110:	sigmoid = 21'b001010101000011110111;
		14'b11110011000111:	sigmoid = 21'b001010101001100101111;
		14'b11110011001000:	sigmoid = 21'b001010101010101100111;
		14'b11110011001001:	sigmoid = 21'b001010101011110100000;
		14'b11110011001010:	sigmoid = 21'b001010101100111011010;
		14'b11110011001011:	sigmoid = 21'b001010101110000010101;
		14'b11110011001100:	sigmoid = 21'b001010101111001010001;
		14'b11110011001101:	sigmoid = 21'b001010110000010001101;
		14'b11110011001110:	sigmoid = 21'b001010110001011001010;
		14'b11110011001111:	sigmoid = 21'b001010110010100001000;
		14'b11110011010000:	sigmoid = 21'b001010110011101000110;
		14'b11110011010001:	sigmoid = 21'b001010110100110000101;
		14'b11110011010010:	sigmoid = 21'b001010110101111000101;
		14'b11110011010011:	sigmoid = 21'b001010110111000000110;
		14'b11110011010100:	sigmoid = 21'b001010111000001001000;
		14'b11110011010101:	sigmoid = 21'b001010111001010001010;
		14'b11110011010110:	sigmoid = 21'b001010111010011001101;
		14'b11110011010111:	sigmoid = 21'b001010111011100010000;
		14'b11110011011000:	sigmoid = 21'b001010111100101010101;
		14'b11110011011001:	sigmoid = 21'b001010111101110011010;
		14'b11110011011010:	sigmoid = 21'b001010111110111100000;
		14'b11110011011011:	sigmoid = 21'b001011000000000100111;
		14'b11110011011100:	sigmoid = 21'b001011000001001101110;
		14'b11110011011101:	sigmoid = 21'b001011000010010110110;
		14'b11110011011110:	sigmoid = 21'b001011000011011111111;
		14'b11110011011111:	sigmoid = 21'b001011000100101001001;
		14'b11110011100000:	sigmoid = 21'b001011000101110010011;
		14'b11110011100001:	sigmoid = 21'b001011000110111011110;
		14'b11110011100010:	sigmoid = 21'b001011001000000101010;
		14'b11110011100011:	sigmoid = 21'b001011001001001110111;
		14'b11110011100100:	sigmoid = 21'b001011001010011000100;
		14'b11110011100101:	sigmoid = 21'b001011001011100010011;
		14'b11110011100110:	sigmoid = 21'b001011001100101100001;
		14'b11110011100111:	sigmoid = 21'b001011001101110110001;
		14'b11110011101000:	sigmoid = 21'b001011001111000000010;
		14'b11110011101001:	sigmoid = 21'b001011010000001010011;
		14'b11110011101010:	sigmoid = 21'b001011010001010100101;
		14'b11110011101011:	sigmoid = 21'b001011010010011110111;
		14'b11110011101100:	sigmoid = 21'b001011010011101001011;
		14'b11110011101101:	sigmoid = 21'b001011010100110011111;
		14'b11110011101110:	sigmoid = 21'b001011010101111110100;
		14'b11110011101111:	sigmoid = 21'b001011010111001001001;
		14'b11110011110000:	sigmoid = 21'b001011011000010100000;
		14'b11110011110001:	sigmoid = 21'b001011011001011110111;
		14'b11110011110010:	sigmoid = 21'b001011011010101001111;
		14'b11110011110011:	sigmoid = 21'b001011011011110101000;
		14'b11110011110100:	sigmoid = 21'b001011011101000000001;
		14'b11110011110101:	sigmoid = 21'b001011011110001011011;
		14'b11110011110110:	sigmoid = 21'b001011011111010110110;
		14'b11110011110111:	sigmoid = 21'b001011100000100010010;
		14'b11110011111000:	sigmoid = 21'b001011100001101101111;
		14'b11110011111001:	sigmoid = 21'b001011100010111001100;
		14'b11110011111010:	sigmoid = 21'b001011100100000101010;
		14'b11110011111011:	sigmoid = 21'b001011100101010001001;
		14'b11110011111100:	sigmoid = 21'b001011100110011101000;
		14'b11110011111101:	sigmoid = 21'b001011100111101001000;
		14'b11110011111110:	sigmoid = 21'b001011101000110101001;
		14'b11110011111111:	sigmoid = 21'b001011101010000001011;
		14'b11110100000000:	sigmoid = 21'b001011101011001101110;
		14'b11110100000001:	sigmoid = 21'b001011101100011010001;
		14'b11110100000010:	sigmoid = 21'b001011101101100110101;
		14'b11110100000011:	sigmoid = 21'b001011101110110011010;
		14'b11110100000100:	sigmoid = 21'b001011101111111111111;
		14'b11110100000101:	sigmoid = 21'b001011110001001100110;
		14'b11110100000110:	sigmoid = 21'b001011110010011001101;
		14'b11110100000111:	sigmoid = 21'b001011110011100110100;
		14'b11110100001000:	sigmoid = 21'b001011110100110011101;
		14'b11110100001001:	sigmoid = 21'b001011110110000000110;
		14'b11110100001010:	sigmoid = 21'b001011110111001110001;
		14'b11110100001011:	sigmoid = 21'b001011111000011011011;
		14'b11110100001100:	sigmoid = 21'b001011111001101000111;
		14'b11110100001101:	sigmoid = 21'b001011111010110110011;
		14'b11110100001110:	sigmoid = 21'b001011111100000100001;
		14'b11110100001111:	sigmoid = 21'b001011111101010001111;
		14'b11110100010000:	sigmoid = 21'b001011111110011111101;
		14'b11110100010001:	sigmoid = 21'b001011111111101101101;
		14'b11110100010010:	sigmoid = 21'b001100000000111011101;
		14'b11110100010011:	sigmoid = 21'b001100000010001001110;
		14'b11110100010100:	sigmoid = 21'b001100000011011000000;
		14'b11110100010101:	sigmoid = 21'b001100000100100110010;
		14'b11110100010110:	sigmoid = 21'b001100000101110100101;
		14'b11110100010111:	sigmoid = 21'b001100000111000011001;
		14'b11110100011000:	sigmoid = 21'b001100001000010001110;
		14'b11110100011001:	sigmoid = 21'b001100001001100000100;
		14'b11110100011010:	sigmoid = 21'b001100001010101111010;
		14'b11110100011011:	sigmoid = 21'b001100001011111110001;
		14'b11110100011100:	sigmoid = 21'b001100001101001101001;
		14'b11110100011101:	sigmoid = 21'b001100001110011100001;
		14'b11110100011110:	sigmoid = 21'b001100001111101011011;
		14'b11110100011111:	sigmoid = 21'b001100010000111010101;
		14'b11110100100000:	sigmoid = 21'b001100010010001010000;
		14'b11110100100001:	sigmoid = 21'b001100010011011001011;
		14'b11110100100010:	sigmoid = 21'b001100010100101001000;
		14'b11110100100011:	sigmoid = 21'b001100010101111000101;
		14'b11110100100100:	sigmoid = 21'b001100010111001000011;
		14'b11110100100101:	sigmoid = 21'b001100011000011000010;
		14'b11110100100110:	sigmoid = 21'b001100011001101000001;
		14'b11110100100111:	sigmoid = 21'b001100011010111000001;
		14'b11110100101000:	sigmoid = 21'b001100011100001000010;
		14'b11110100101001:	sigmoid = 21'b001100011101011000100;
		14'b11110100101010:	sigmoid = 21'b001100011110101000111;
		14'b11110100101011:	sigmoid = 21'b001100011111111001010;
		14'b11110100101100:	sigmoid = 21'b001100100001001001110;
		14'b11110100101101:	sigmoid = 21'b001100100010011010011;
		14'b11110100101110:	sigmoid = 21'b001100100011101011000;
		14'b11110100101111:	sigmoid = 21'b001100100100111011111;
		14'b11110100110000:	sigmoid = 21'b001100100110001100110;
		14'b11110100110001:	sigmoid = 21'b001100100111011101110;
		14'b11110100110010:	sigmoid = 21'b001100101000101110111;
		14'b11110100110011:	sigmoid = 21'b001100101010000000000;
		14'b11110100110100:	sigmoid = 21'b001100101011010001010;
		14'b11110100110101:	sigmoid = 21'b001100101100100010101;
		14'b11110100110110:	sigmoid = 21'b001100101101110100001;
		14'b11110100110111:	sigmoid = 21'b001100101111000101101;
		14'b11110100111000:	sigmoid = 21'b001100110000010111011;
		14'b11110100111001:	sigmoid = 21'b001100110001101001001;
		14'b11110100111010:	sigmoid = 21'b001100110010111011000;
		14'b11110100111011:	sigmoid = 21'b001100110100001100111;
		14'b11110100111100:	sigmoid = 21'b001100110101011110111;
		14'b11110100111101:	sigmoid = 21'b001100110110110001001;
		14'b11110100111110:	sigmoid = 21'b001100111000000011010;
		14'b11110100111111:	sigmoid = 21'b001100111001010101101;
		14'b11110101000000:	sigmoid = 21'b001100111010101000001;
		14'b11110101000001:	sigmoid = 21'b001100111011111010101;
		14'b11110101000010:	sigmoid = 21'b001100111101001101010;
		14'b11110101000011:	sigmoid = 21'b001100111110011111111;
		14'b11110101000100:	sigmoid = 21'b001100111111110010110;
		14'b11110101000101:	sigmoid = 21'b001101000001000101101;
		14'b11110101000110:	sigmoid = 21'b001101000010011000101;
		14'b11110101000111:	sigmoid = 21'b001101000011101011110;
		14'b11110101001000:	sigmoid = 21'b001101000100111111000;
		14'b11110101001001:	sigmoid = 21'b001101000110010010010;
		14'b11110101001010:	sigmoid = 21'b001101000111100101101;
		14'b11110101001011:	sigmoid = 21'b001101001000111001001;
		14'b11110101001100:	sigmoid = 21'b001101001010001100101;
		14'b11110101001101:	sigmoid = 21'b001101001011100000011;
		14'b11110101001110:	sigmoid = 21'b001101001100110100001;
		14'b11110101001111:	sigmoid = 21'b001101001110001000000;
		14'b11110101010000:	sigmoid = 21'b001101001111011100000;
		14'b11110101010001:	sigmoid = 21'b001101010000110000000;
		14'b11110101010010:	sigmoid = 21'b001101010010000100010;
		14'b11110101010011:	sigmoid = 21'b001101010011011000100;
		14'b11110101010100:	sigmoid = 21'b001101010100101100110;
		14'b11110101010101:	sigmoid = 21'b001101010110000001010;
		14'b11110101010110:	sigmoid = 21'b001101010111010101110;
		14'b11110101010111:	sigmoid = 21'b001101011000101010011;
		14'b11110101011000:	sigmoid = 21'b001101011001111111001;
		14'b11110101011001:	sigmoid = 21'b001101011011010100000;
		14'b11110101011010:	sigmoid = 21'b001101011100101000111;
		14'b11110101011011:	sigmoid = 21'b001101011101111110000;
		14'b11110101011100:	sigmoid = 21'b001101011111010011000;
		14'b11110101011101:	sigmoid = 21'b001101100000101000010;
		14'b11110101011110:	sigmoid = 21'b001101100001111101101;
		14'b11110101011111:	sigmoid = 21'b001101100011010011000;
		14'b11110101100000:	sigmoid = 21'b001101100100101000100;
		14'b11110101100001:	sigmoid = 21'b001101100101111110001;
		14'b11110101100010:	sigmoid = 21'b001101100111010011110;
		14'b11110101100011:	sigmoid = 21'b001101101000101001101;
		14'b11110101100100:	sigmoid = 21'b001101101001111111100;
		14'b11110101100101:	sigmoid = 21'b001101101011010101100;
		14'b11110101100110:	sigmoid = 21'b001101101100101011100;
		14'b11110101100111:	sigmoid = 21'b001101101110000001110;
		14'b11110101101000:	sigmoid = 21'b001101101111011000000;
		14'b11110101101001:	sigmoid = 21'b001101110000101110011;
		14'b11110101101010:	sigmoid = 21'b001101110010000100111;
		14'b11110101101011:	sigmoid = 21'b001101110011011011011;
		14'b11110101101100:	sigmoid = 21'b001101110100110010001;
		14'b11110101101101:	sigmoid = 21'b001101110110001000111;
		14'b11110101101110:	sigmoid = 21'b001101110111011111101;
		14'b11110101101111:	sigmoid = 21'b001101111000110110101;
		14'b11110101110000:	sigmoid = 21'b001101111010001101101;
		14'b11110101110001:	sigmoid = 21'b001101111011100100110;
		14'b11110101110010:	sigmoid = 21'b001101111100111100000;
		14'b11110101110011:	sigmoid = 21'b001101111110010011011;
		14'b11110101110100:	sigmoid = 21'b001101111111101010110;
		14'b11110101110101:	sigmoid = 21'b001110000001000010011;
		14'b11110101110110:	sigmoid = 21'b001110000010011010000;
		14'b11110101110111:	sigmoid = 21'b001110000011110001101;
		14'b11110101111000:	sigmoid = 21'b001110000101001001100;
		14'b11110101111001:	sigmoid = 21'b001110000110100001011;
		14'b11110101111010:	sigmoid = 21'b001110000111111001011;
		14'b11110101111011:	sigmoid = 21'b001110001001010001100;
		14'b11110101111100:	sigmoid = 21'b001110001010101001110;
		14'b11110101111101:	sigmoid = 21'b001110001100000010000;
		14'b11110101111110:	sigmoid = 21'b001110001101011010011;
		14'b11110101111111:	sigmoid = 21'b001110001110110010111;
		14'b11110110000000:	sigmoid = 21'b001110010000001011100;
		14'b11110110000001:	sigmoid = 21'b001110010001100100001;
		14'b11110110000010:	sigmoid = 21'b001110010010111100111;
		14'b11110110000011:	sigmoid = 21'b001110010100010101110;
		14'b11110110000100:	sigmoid = 21'b001110010101101110110;
		14'b11110110000101:	sigmoid = 21'b001110010111000111110;
		14'b11110110000110:	sigmoid = 21'b001110011000100001000;
		14'b11110110000111:	sigmoid = 21'b001110011001111010010;
		14'b11110110001000:	sigmoid = 21'b001110011011010011100;
		14'b11110110001001:	sigmoid = 21'b001110011100101101000;
		14'b11110110001010:	sigmoid = 21'b001110011110000110100;
		14'b11110110001011:	sigmoid = 21'b001110011111100000001;
		14'b11110110001100:	sigmoid = 21'b001110100000111001111;
		14'b11110110001101:	sigmoid = 21'b001110100010010011110;
		14'b11110110001110:	sigmoid = 21'b001110100011101101101;
		14'b11110110001111:	sigmoid = 21'b001110100101000111101;
		14'b11110110010000:	sigmoid = 21'b001110100110100001110;
		14'b11110110010001:	sigmoid = 21'b001110100111111100000;
		14'b11110110010010:	sigmoid = 21'b001110101001010110011;
		14'b11110110010011:	sigmoid = 21'b001110101010110000110;
		14'b11110110010100:	sigmoid = 21'b001110101100001011010;
		14'b11110110010101:	sigmoid = 21'b001110101101100101110;
		14'b11110110010110:	sigmoid = 21'b001110101111000000100;
		14'b11110110010111:	sigmoid = 21'b001110110000011011010;
		14'b11110110011000:	sigmoid = 21'b001110110001110110001;
		14'b11110110011001:	sigmoid = 21'b001110110011010001001;
		14'b11110110011010:	sigmoid = 21'b001110110100101100010;
		14'b11110110011011:	sigmoid = 21'b001110110110000111011;
		14'b11110110011100:	sigmoid = 21'b001110110111100010101;
		14'b11110110011101:	sigmoid = 21'b001110111000111110000;
		14'b11110110011110:	sigmoid = 21'b001110111010011001100;
		14'b11110110011111:	sigmoid = 21'b001110111011110101000;
		14'b11110110100000:	sigmoid = 21'b001110111101010000101;
		14'b11110110100001:	sigmoid = 21'b001110111110101100011;
		14'b11110110100010:	sigmoid = 21'b001111000000001000010;
		14'b11110110100011:	sigmoid = 21'b001111000001100100001;
		14'b11110110100100:	sigmoid = 21'b001111000011000000010;
		14'b11110110100101:	sigmoid = 21'b001111000100011100011;
		14'b11110110100110:	sigmoid = 21'b001111000101111000100;
		14'b11110110100111:	sigmoid = 21'b001111000111010100111;
		14'b11110110101000:	sigmoid = 21'b001111001000110001010;
		14'b11110110101001:	sigmoid = 21'b001111001010001101110;
		14'b11110110101010:	sigmoid = 21'b001111001011101010011;
		14'b11110110101011:	sigmoid = 21'b001111001101000111000;
		14'b11110110101100:	sigmoid = 21'b001111001110100011111;
		14'b11110110101101:	sigmoid = 21'b001111010000000000110;
		14'b11110110101110:	sigmoid = 21'b001111010001011101110;
		14'b11110110101111:	sigmoid = 21'b001111010010111010110;
		14'b11110110110000:	sigmoid = 21'b001111010100010111111;
		14'b11110110110001:	sigmoid = 21'b001111010101110101010;
		14'b11110110110010:	sigmoid = 21'b001111010111010010100;
		14'b11110110110011:	sigmoid = 21'b001111011000110000000;
		14'b11110110110100:	sigmoid = 21'b001111011010001101100;
		14'b11110110110101:	sigmoid = 21'b001111011011101011010;
		14'b11110110110110:	sigmoid = 21'b001111011101001000111;
		14'b11110110110111:	sigmoid = 21'b001111011110100110110;
		14'b11110110111000:	sigmoid = 21'b001111100000000100110;
		14'b11110110111001:	sigmoid = 21'b001111100001100010110;
		14'b11110110111010:	sigmoid = 21'b001111100011000000111;
		14'b11110110111011:	sigmoid = 21'b001111100100011111000;
		14'b11110110111100:	sigmoid = 21'b001111100101111101011;
		14'b11110110111101:	sigmoid = 21'b001111100111011011110;
		14'b11110110111110:	sigmoid = 21'b001111101000111010010;
		14'b11110110111111:	sigmoid = 21'b001111101010011000111;
		14'b11110111000000:	sigmoid = 21'b001111101011110111100;
		14'b11110111000001:	sigmoid = 21'b001111101101010110010;
		14'b11110111000010:	sigmoid = 21'b001111101110110101001;
		14'b11110111000011:	sigmoid = 21'b001111110000010100001;
		14'b11110111000100:	sigmoid = 21'b001111110001110011001;
		14'b11110111000101:	sigmoid = 21'b001111110011010010011;
		14'b11110111000110:	sigmoid = 21'b001111110100110001101;
		14'b11110111000111:	sigmoid = 21'b001111110110010000111;
		14'b11110111001000:	sigmoid = 21'b001111110111110000011;
		14'b11110111001001:	sigmoid = 21'b001111111001001111111;
		14'b11110111001010:	sigmoid = 21'b001111111010101111100;
		14'b11110111001011:	sigmoid = 21'b001111111100001111010;
		14'b11110111001100:	sigmoid = 21'b001111111101101111000;
		14'b11110111001101:	sigmoid = 21'b001111111111001111000;
		14'b11110111001110:	sigmoid = 21'b010000000000101111000;
		14'b11110111001111:	sigmoid = 21'b010000000010001111000;
		14'b11110111010000:	sigmoid = 21'b010000000011101111010;
		14'b11110111010001:	sigmoid = 21'b010000000101001111100;
		14'b11110111010010:	sigmoid = 21'b010000000110101111111;
		14'b11110111010011:	sigmoid = 21'b010000001000010000011;
		14'b11110111010100:	sigmoid = 21'b010000001001110000111;
		14'b11110111010101:	sigmoid = 21'b010000001011010001100;
		14'b11110111010110:	sigmoid = 21'b010000001100110010010;
		14'b11110111010111:	sigmoid = 21'b010000001110010011001;
		14'b11110111011000:	sigmoid = 21'b010000001111110100001;
		14'b11110111011001:	sigmoid = 21'b010000010001010101001;
		14'b11110111011010:	sigmoid = 21'b010000010010110110010;
		14'b11110111011011:	sigmoid = 21'b010000010100010111100;
		14'b11110111011100:	sigmoid = 21'b010000010101111000110;
		14'b11110111011101:	sigmoid = 21'b010000010111011010001;
		14'b11110111011110:	sigmoid = 21'b010000011000111011101;
		14'b11110111011111:	sigmoid = 21'b010000011010011101010;
		14'b11110111100000:	sigmoid = 21'b010000011011111110111;
		14'b11110111100001:	sigmoid = 21'b010000011101100000101;
		14'b11110111100010:	sigmoid = 21'b010000011111000010100;
		14'b11110111100011:	sigmoid = 21'b010000100000100100100;
		14'b11110111100100:	sigmoid = 21'b010000100010000110100;
		14'b11110111100101:	sigmoid = 21'b010000100011101000110;
		14'b11110111100110:	sigmoid = 21'b010000100101001010111;
		14'b11110111100111:	sigmoid = 21'b010000100110101101010;
		14'b11110111101000:	sigmoid = 21'b010000101000001111101;
		14'b11110111101001:	sigmoid = 21'b010000101001110010001;
		14'b11110111101010:	sigmoid = 21'b010000101011010100110;
		14'b11110111101011:	sigmoid = 21'b010000101100110111100;
		14'b11110111101100:	sigmoid = 21'b010000101110011010010;
		14'b11110111101101:	sigmoid = 21'b010000101111111101001;
		14'b11110111101110:	sigmoid = 21'b010000110001100000001;
		14'b11110111101111:	sigmoid = 21'b010000110011000011010;
		14'b11110111110000:	sigmoid = 21'b010000110100100110011;
		14'b11110111110001:	sigmoid = 21'b010000110110001001101;
		14'b11110111110010:	sigmoid = 21'b010000110111101101000;
		14'b11110111110011:	sigmoid = 21'b010000111001010000011;
		14'b11110111110100:	sigmoid = 21'b010000111010110011111;
		14'b11110111110101:	sigmoid = 21'b010000111100010111100;
		14'b11110111110110:	sigmoid = 21'b010000111101111011010;
		14'b11110111110111:	sigmoid = 21'b010000111111011111000;
		14'b11110111111000:	sigmoid = 21'b010001000001000010111;
		14'b11110111111001:	sigmoid = 21'b010001000010100110111;
		14'b11110111111010:	sigmoid = 21'b010001000100001011000;
		14'b11110111111011:	sigmoid = 21'b010001000101101111001;
		14'b11110111111100:	sigmoid = 21'b010001000111010011011;
		14'b11110111111101:	sigmoid = 21'b010001001000110111110;
		14'b11110111111110:	sigmoid = 21'b010001001010011100001;
		14'b11110111111111:	sigmoid = 21'b010001001100000000110;
		14'b11111000000000:	sigmoid = 21'b010001001101100101011;
		14'b11111000000001:	sigmoid = 21'b010001001111001010000;
		14'b11111000000010:	sigmoid = 21'b010001010000101110111;
		14'b11111000000011:	sigmoid = 21'b010001010010010011110;
		14'b11111000000100:	sigmoid = 21'b010001010011111000110;
		14'b11111000000101:	sigmoid = 21'b010001010101011101110;
		14'b11111000000110:	sigmoid = 21'b010001010111000011000;
		14'b11111000000111:	sigmoid = 21'b010001011000101000010;
		14'b11111000001000:	sigmoid = 21'b010001011010001101100;
		14'b11111000001001:	sigmoid = 21'b010001011011110011000;
		14'b11111000001010:	sigmoid = 21'b010001011101011000100;
		14'b11111000001011:	sigmoid = 21'b010001011110111110001;
		14'b11111000001100:	sigmoid = 21'b010001100000100011111;
		14'b11111000001101:	sigmoid = 21'b010001100010001001101;
		14'b11111000001110:	sigmoid = 21'b010001100011101111100;
		14'b11111000001111:	sigmoid = 21'b010001100101010101100;
		14'b11111000010000:	sigmoid = 21'b010001100110111011100;
		14'b11111000010001:	sigmoid = 21'b010001101000100001110;
		14'b11111000010010:	sigmoid = 21'b010001101010001000000;
		14'b11111000010011:	sigmoid = 21'b010001101011101110010;
		14'b11111000010100:	sigmoid = 21'b010001101101010100110;
		14'b11111000010101:	sigmoid = 21'b010001101110111011010;
		14'b11111000010110:	sigmoid = 21'b010001110000100001111;
		14'b11111000010111:	sigmoid = 21'b010001110010001000100;
		14'b11111000011000:	sigmoid = 21'b010001110011101111010;
		14'b11111000011001:	sigmoid = 21'b010001110101010110001;
		14'b11111000011010:	sigmoid = 21'b010001110110111101001;
		14'b11111000011011:	sigmoid = 21'b010001111000100100001;
		14'b11111000011100:	sigmoid = 21'b010001111010001011010;
		14'b11111000011101:	sigmoid = 21'b010001111011110010100;
		14'b11111000011110:	sigmoid = 21'b010001111101011001111;
		14'b11111000011111:	sigmoid = 21'b010001111111000001010;
		14'b11111000100000:	sigmoid = 21'b010010000000101000110;
		14'b11111000100001:	sigmoid = 21'b010010000010010000010;
		14'b11111000100010:	sigmoid = 21'b010010000011111000000;
		14'b11111000100011:	sigmoid = 21'b010010000101011111110;
		14'b11111000100100:	sigmoid = 21'b010010000111000111101;
		14'b11111000100101:	sigmoid = 21'b010010001000101111100;
		14'b11111000100110:	sigmoid = 21'b010010001010010111100;
		14'b11111000100111:	sigmoid = 21'b010010001011111111101;
		14'b11111000101000:	sigmoid = 21'b010010001101100111111;
		14'b11111000101001:	sigmoid = 21'b010010001111010000001;
		14'b11111000101010:	sigmoid = 21'b010010010000111000100;
		14'b11111000101011:	sigmoid = 21'b010010010010100001000;
		14'b11111000101100:	sigmoid = 21'b010010010100001001100;
		14'b11111000101101:	sigmoid = 21'b010010010101110010001;
		14'b11111000101110:	sigmoid = 21'b010010010111011010111;
		14'b11111000101111:	sigmoid = 21'b010010011001000011101;
		14'b11111000110000:	sigmoid = 21'b010010011010101100100;
		14'b11111000110001:	sigmoid = 21'b010010011100010101100;
		14'b11111000110010:	sigmoid = 21'b010010011101111110101;
		14'b11111000110011:	sigmoid = 21'b010010011111100111110;
		14'b11111000110100:	sigmoid = 21'b010010100001010001000;
		14'b11111000110101:	sigmoid = 21'b010010100010111010011;
		14'b11111000110110:	sigmoid = 21'b010010100100100011110;
		14'b11111000110111:	sigmoid = 21'b010010100110001101010;
		14'b11111000111000:	sigmoid = 21'b010010100111110110111;
		14'b11111000111001:	sigmoid = 21'b010010101001100000100;
		14'b11111000111010:	sigmoid = 21'b010010101011001010010;
		14'b11111000111011:	sigmoid = 21'b010010101100110100001;
		14'b11111000111100:	sigmoid = 21'b010010101110011110000;
		14'b11111000111101:	sigmoid = 21'b010010110000001000000;
		14'b11111000111110:	sigmoid = 21'b010010110001110010001;
		14'b11111000111111:	sigmoid = 21'b010010110011011100011;
		14'b11111001000000:	sigmoid = 21'b010010110101000110101;
		14'b11111001000001:	sigmoid = 21'b010010110110110001000;
		14'b11111001000010:	sigmoid = 21'b010010111000011011011;
		14'b11111001000011:	sigmoid = 21'b010010111010000110000;
		14'b11111001000100:	sigmoid = 21'b010010111011110000101;
		14'b11111001000101:	sigmoid = 21'b010010111101011011010;
		14'b11111001000110:	sigmoid = 21'b010010111111000110001;
		14'b11111001000111:	sigmoid = 21'b010011000000110001000;
		14'b11111001001000:	sigmoid = 21'b010011000010011011111;
		14'b11111001001001:	sigmoid = 21'b010011000100000111000;
		14'b11111001001010:	sigmoid = 21'b010011000101110010001;
		14'b11111001001011:	sigmoid = 21'b010011000111011101010;
		14'b11111001001100:	sigmoid = 21'b010011001001001000101;
		14'b11111001001101:	sigmoid = 21'b010011001010110100000;
		14'b11111001001110:	sigmoid = 21'b010011001100011111011;
		14'b11111001001111:	sigmoid = 21'b010011001110001011000;
		14'b11111001010000:	sigmoid = 21'b010011001111110110101;
		14'b11111001010001:	sigmoid = 21'b010011010001100010010;
		14'b11111001010010:	sigmoid = 21'b010011010011001110001;
		14'b11111001010011:	sigmoid = 21'b010011010100111010000;
		14'b11111001010100:	sigmoid = 21'b010011010110100110000;
		14'b11111001010101:	sigmoid = 21'b010011011000010010000;
		14'b11111001010110:	sigmoid = 21'b010011011001111110001;
		14'b11111001010111:	sigmoid = 21'b010011011011101010011;
		14'b11111001011000:	sigmoid = 21'b010011011101010110101;
		14'b11111001011001:	sigmoid = 21'b010011011111000011000;
		14'b11111001011010:	sigmoid = 21'b010011100000101111100;
		14'b11111001011011:	sigmoid = 21'b010011100010011100000;
		14'b11111001011100:	sigmoid = 21'b010011100100001000101;
		14'b11111001011101:	sigmoid = 21'b010011100101110101011;
		14'b11111001011110:	sigmoid = 21'b010011100111100010001;
		14'b11111001011111:	sigmoid = 21'b010011101001001111000;
		14'b11111001100000:	sigmoid = 21'b010011101010111100000;
		14'b11111001100001:	sigmoid = 21'b010011101100101001000;
		14'b11111001100010:	sigmoid = 21'b010011101110010110001;
		14'b11111001100011:	sigmoid = 21'b010011110000000011011;
		14'b11111001100100:	sigmoid = 21'b010011110001110000101;
		14'b11111001100101:	sigmoid = 21'b010011110011011110000;
		14'b11111001100110:	sigmoid = 21'b010011110101001011100;
		14'b11111001100111:	sigmoid = 21'b010011110110111001000;
		14'b11111001101000:	sigmoid = 21'b010011111000100110101;
		14'b11111001101001:	sigmoid = 21'b010011111010010100010;
		14'b11111001101010:	sigmoid = 21'b010011111100000010001;
		14'b11111001101011:	sigmoid = 21'b010011111101101111111;
		14'b11111001101100:	sigmoid = 21'b010011111111011101111;
		14'b11111001101101:	sigmoid = 21'b010100000001001011111;
		14'b11111001101110:	sigmoid = 21'b010100000010111010000;
		14'b11111001101111:	sigmoid = 21'b010100000100101000001;
		14'b11111001110000:	sigmoid = 21'b010100000110010110011;
		14'b11111001110001:	sigmoid = 21'b010100001000000100110;
		14'b11111001110010:	sigmoid = 21'b010100001001110011001;
		14'b11111001110011:	sigmoid = 21'b010100001011100001101;
		14'b11111001110100:	sigmoid = 21'b010100001101010000010;
		14'b11111001110101:	sigmoid = 21'b010100001110111110111;
		14'b11111001110110:	sigmoid = 21'b010100010000101101101;
		14'b11111001110111:	sigmoid = 21'b010100010010011100011;
		14'b11111001111000:	sigmoid = 21'b010100010100001011011;
		14'b11111001111001:	sigmoid = 21'b010100010101111010010;
		14'b11111001111010:	sigmoid = 21'b010100010111101001011;
		14'b11111001111011:	sigmoid = 21'b010100011001011000100;
		14'b11111001111100:	sigmoid = 21'b010100011011000111110;
		14'b11111001111101:	sigmoid = 21'b010100011100110111000;
		14'b11111001111110:	sigmoid = 21'b010100011110100110011;
		14'b11111001111111:	sigmoid = 21'b010100100000010101110;
		14'b11111010000000:	sigmoid = 21'b010100100010000101011;
		14'b11111010000001:	sigmoid = 21'b010100100011110100111;
		14'b11111010000010:	sigmoid = 21'b010100100101100100101;
		14'b11111010000011:	sigmoid = 21'b010100100111010100011;
		14'b11111010000100:	sigmoid = 21'b010100101001000100010;
		14'b11111010000101:	sigmoid = 21'b010100101010110100001;
		14'b11111010000110:	sigmoid = 21'b010100101100100100001;
		14'b11111010000111:	sigmoid = 21'b010100101110010100001;
		14'b11111010001000:	sigmoid = 21'b010100110000000100010;
		14'b11111010001001:	sigmoid = 21'b010100110001110100100;
		14'b11111010001010:	sigmoid = 21'b010100110011100100111;
		14'b11111010001011:	sigmoid = 21'b010100110101010101010;
		14'b11111010001100:	sigmoid = 21'b010100110111000101101;
		14'b11111010001101:	sigmoid = 21'b010100111000110110001;
		14'b11111010001110:	sigmoid = 21'b010100111010100110110;
		14'b11111010001111:	sigmoid = 21'b010100111100010111100;
		14'b11111010010000:	sigmoid = 21'b010100111110001000010;
		14'b11111010010001:	sigmoid = 21'b010100111111111001000;
		14'b11111010010010:	sigmoid = 21'b010101000001101010000;
		14'b11111010010011:	sigmoid = 21'b010101000011011011000;
		14'b11111010010100:	sigmoid = 21'b010101000101001100000;
		14'b11111010010101:	sigmoid = 21'b010101000110111101001;
		14'b11111010010110:	sigmoid = 21'b010101001000101110011;
		14'b11111010010111:	sigmoid = 21'b010101001010011111101;
		14'b11111010011000:	sigmoid = 21'b010101001100010001000;
		14'b11111010011001:	sigmoid = 21'b010101001110000010011;
		14'b11111010011010:	sigmoid = 21'b010101001111110011111;
		14'b11111010011011:	sigmoid = 21'b010101010001100101100;
		14'b11111010011100:	sigmoid = 21'b010101010011010111001;
		14'b11111010011101:	sigmoid = 21'b010101010101001000111;
		14'b11111010011110:	sigmoid = 21'b010101010110111010110;
		14'b11111010011111:	sigmoid = 21'b010101011000101100101;
		14'b11111010100000:	sigmoid = 21'b010101011010011110100;
		14'b11111010100001:	sigmoid = 21'b010101011100010000101;
		14'b11111010100010:	sigmoid = 21'b010101011110000010101;
		14'b11111010100011:	sigmoid = 21'b010101011111110100111;
		14'b11111010100100:	sigmoid = 21'b010101100001100111001;
		14'b11111010100101:	sigmoid = 21'b010101100011011001011;
		14'b11111010100110:	sigmoid = 21'b010101100101001011111;
		14'b11111010100111:	sigmoid = 21'b010101100110111110010;
		14'b11111010101000:	sigmoid = 21'b010101101000110000111;
		14'b11111010101001:	sigmoid = 21'b010101101010100011100;
		14'b11111010101010:	sigmoid = 21'b010101101100010110001;
		14'b11111010101011:	sigmoid = 21'b010101101110001000111;
		14'b11111010101100:	sigmoid = 21'b010101101111111011110;
		14'b11111010101101:	sigmoid = 21'b010101110001101110101;
		14'b11111010101110:	sigmoid = 21'b010101110011100001101;
		14'b11111010101111:	sigmoid = 21'b010101110101010100101;
		14'b11111010110000:	sigmoid = 21'b010101110111000111110;
		14'b11111010110001:	sigmoid = 21'b010101111000111010111;
		14'b11111010110010:	sigmoid = 21'b010101111010101110001;
		14'b11111010110011:	sigmoid = 21'b010101111100100001100;
		14'b11111010110100:	sigmoid = 21'b010101111110010100111;
		14'b11111010110101:	sigmoid = 21'b010110000000001000011;
		14'b11111010110110:	sigmoid = 21'b010110000001111011111;
		14'b11111010110111:	sigmoid = 21'b010110000011101111100;
		14'b11111010111000:	sigmoid = 21'b010110000101100011010;
		14'b11111010111001:	sigmoid = 21'b010110000111010111000;
		14'b11111010111010:	sigmoid = 21'b010110001001001010110;
		14'b11111010111011:	sigmoid = 21'b010110001010111110101;
		14'b11111010111100:	sigmoid = 21'b010110001100110010101;
		14'b11111010111101:	sigmoid = 21'b010110001110100110101;
		14'b11111010111110:	sigmoid = 21'b010110010000011010110;
		14'b11111010111111:	sigmoid = 21'b010110010010001110111;
		14'b11111011000000:	sigmoid = 21'b010110010100000011001;
		14'b11111011000001:	sigmoid = 21'b010110010101110111100;
		14'b11111011000010:	sigmoid = 21'b010110010111101011111;
		14'b11111011000011:	sigmoid = 21'b010110011001100000010;
		14'b11111011000100:	sigmoid = 21'b010110011011010100110;
		14'b11111011000101:	sigmoid = 21'b010110011101001001011;
		14'b11111011000110:	sigmoid = 21'b010110011110111110000;
		14'b11111011000111:	sigmoid = 21'b010110100000110010110;
		14'b11111011001000:	sigmoid = 21'b010110100010100111100;
		14'b11111011001001:	sigmoid = 21'b010110100100011100011;
		14'b11111011001010:	sigmoid = 21'b010110100110010001010;
		14'b11111011001011:	sigmoid = 21'b010110101000000110010;
		14'b11111011001100:	sigmoid = 21'b010110101001111011011;
		14'b11111011001101:	sigmoid = 21'b010110101011110000100;
		14'b11111011001110:	sigmoid = 21'b010110101101100101101;
		14'b11111011001111:	sigmoid = 21'b010110101111011010111;
		14'b11111011010000:	sigmoid = 21'b010110110001010000010;
		14'b11111011010001:	sigmoid = 21'b010110110011000101101;
		14'b11111011010010:	sigmoid = 21'b010110110100111011000;
		14'b11111011010011:	sigmoid = 21'b010110110110110000100;
		14'b11111011010100:	sigmoid = 21'b010110111000100110001;
		14'b11111011010101:	sigmoid = 21'b010110111010011011110;
		14'b11111011010110:	sigmoid = 21'b010110111100010001100;
		14'b11111011010111:	sigmoid = 21'b010110111110000111010;
		14'b11111011011000:	sigmoid = 21'b010110111111111101001;
		14'b11111011011001:	sigmoid = 21'b010111000001110011000;
		14'b11111011011010:	sigmoid = 21'b010111000011101001000;
		14'b11111011011011:	sigmoid = 21'b010111000101011111000;
		14'b11111011011100:	sigmoid = 21'b010111000111010101001;
		14'b11111011011101:	sigmoid = 21'b010111001001001011010;
		14'b11111011011110:	sigmoid = 21'b010111001011000001100;
		14'b11111011011111:	sigmoid = 21'b010111001100110111110;
		14'b11111011100000:	sigmoid = 21'b010111001110101110001;
		14'b11111011100001:	sigmoid = 21'b010111010000100100100;
		14'b11111011100010:	sigmoid = 21'b010111010010011011000;
		14'b11111011100011:	sigmoid = 21'b010111010100010001101;
		14'b11111011100100:	sigmoid = 21'b010111010110001000001;
		14'b11111011100101:	sigmoid = 21'b010111010111111110111;
		14'b11111011100110:	sigmoid = 21'b010111011001110101101;
		14'b11111011100111:	sigmoid = 21'b010111011011101100011;
		14'b11111011101000:	sigmoid = 21'b010111011101100011010;
		14'b11111011101001:	sigmoid = 21'b010111011111011010001;
		14'b11111011101010:	sigmoid = 21'b010111100001010001001;
		14'b11111011101011:	sigmoid = 21'b010111100011001000001;
		14'b11111011101100:	sigmoid = 21'b010111100100111111010;
		14'b11111011101101:	sigmoid = 21'b010111100110110110100;
		14'b11111011101110:	sigmoid = 21'b010111101000101101101;
		14'b11111011101111:	sigmoid = 21'b010111101010100101000;
		14'b11111011110000:	sigmoid = 21'b010111101100011100010;
		14'b11111011110001:	sigmoid = 21'b010111101110010011110;
		14'b11111011110010:	sigmoid = 21'b010111110000001011001;
		14'b11111011110011:	sigmoid = 21'b010111110010000010110;
		14'b11111011110100:	sigmoid = 21'b010111110011111010010;
		14'b11111011110101:	sigmoid = 21'b010111110101110010000;
		14'b11111011110110:	sigmoid = 21'b010111110111101001101;
		14'b11111011110111:	sigmoid = 21'b010111111001100001011;
		14'b11111011111000:	sigmoid = 21'b010111111011011001010;
		14'b11111011111001:	sigmoid = 21'b010111111101010001001;
		14'b11111011111010:	sigmoid = 21'b010111111111001001001;
		14'b11111011111011:	sigmoid = 21'b011000000001000001001;
		14'b11111011111100:	sigmoid = 21'b011000000010111001001;
		14'b11111011111101:	sigmoid = 21'b011000000100110001010;
		14'b11111011111110:	sigmoid = 21'b011000000110101001011;
		14'b11111011111111:	sigmoid = 21'b011000001000100001101;
		14'b11111100000000:	sigmoid = 21'b011000001010011010000;
		14'b11111100000001:	sigmoid = 21'b011000001100010010010;
		14'b11111100000010:	sigmoid = 21'b011000001110001010110;
		14'b11111100000011:	sigmoid = 21'b011000010000000011001;
		14'b11111100000100:	sigmoid = 21'b011000010001111011110;
		14'b11111100000101:	sigmoid = 21'b011000010011110100010;
		14'b11111100000110:	sigmoid = 21'b011000010101101100111;
		14'b11111100000111:	sigmoid = 21'b011000010111100101101;
		14'b11111100001000:	sigmoid = 21'b011000011001011110011;
		14'b11111100001001:	sigmoid = 21'b011000011011010111001;
		14'b11111100001010:	sigmoid = 21'b011000011101010000000;
		14'b11111100001011:	sigmoid = 21'b011000011111001001000;
		14'b11111100001100:	sigmoid = 21'b011000100001000001111;
		14'b11111100001101:	sigmoid = 21'b011000100010111010111;
		14'b11111100001110:	sigmoid = 21'b011000100100110100000;
		14'b11111100001111:	sigmoid = 21'b011000100110101101001;
		14'b11111100010000:	sigmoid = 21'b011000101000100110011;
		14'b11111100010001:	sigmoid = 21'b011000101010011111101;
		14'b11111100010010:	sigmoid = 21'b011000101100011000111;
		14'b11111100010011:	sigmoid = 21'b011000101110010010010;
		14'b11111100010100:	sigmoid = 21'b011000110000001011101;
		14'b11111100010101:	sigmoid = 21'b011000110010000101001;
		14'b11111100010110:	sigmoid = 21'b011000110011111110101;
		14'b11111100010111:	sigmoid = 21'b011000110101111000010;
		14'b11111100011000:	sigmoid = 21'b011000110111110001111;
		14'b11111100011001:	sigmoid = 21'b011000111001101011100;
		14'b11111100011010:	sigmoid = 21'b011000111011100101010;
		14'b11111100011011:	sigmoid = 21'b011000111101011111000;
		14'b11111100011100:	sigmoid = 21'b011000111111011000111;
		14'b11111100011101:	sigmoid = 21'b011001000001010010110;
		14'b11111100011110:	sigmoid = 21'b011001000011001100101;
		14'b11111100011111:	sigmoid = 21'b011001000101000110101;
		14'b11111100100000:	sigmoid = 21'b011001000111000000101;
		14'b11111100100001:	sigmoid = 21'b011001001000111010110;
		14'b11111100100010:	sigmoid = 21'b011001001010110100111;
		14'b11111100100011:	sigmoid = 21'b011001001100101111001;
		14'b11111100100100:	sigmoid = 21'b011001001110101001011;
		14'b11111100100101:	sigmoid = 21'b011001010000100011101;
		14'b11111100100110:	sigmoid = 21'b011001010010011110000;
		14'b11111100100111:	sigmoid = 21'b011001010100011000011;
		14'b11111100101000:	sigmoid = 21'b011001010110010010111;
		14'b11111100101001:	sigmoid = 21'b011001011000001101011;
		14'b11111100101010:	sigmoid = 21'b011001011010000111111;
		14'b11111100101011:	sigmoid = 21'b011001011100000010100;
		14'b11111100101100:	sigmoid = 21'b011001011101111101001;
		14'b11111100101101:	sigmoid = 21'b011001011111110111110;
		14'b11111100101110:	sigmoid = 21'b011001100001110010100;
		14'b11111100101111:	sigmoid = 21'b011001100011101101011;
		14'b11111100110000:	sigmoid = 21'b011001100101101000001;
		14'b11111100110001:	sigmoid = 21'b011001100111100011000;
		14'b11111100110010:	sigmoid = 21'b011001101001011110000;
		14'b11111100110011:	sigmoid = 21'b011001101011011001000;
		14'b11111100110100:	sigmoid = 21'b011001101101010100000;
		14'b11111100110101:	sigmoid = 21'b011001101111001111000;
		14'b11111100110110:	sigmoid = 21'b011001110001001010001;
		14'b11111100110111:	sigmoid = 21'b011001110011000101011;
		14'b11111100111000:	sigmoid = 21'b011001110101000000101;
		14'b11111100111001:	sigmoid = 21'b011001110110111011111;
		14'b11111100111010:	sigmoid = 21'b011001111000110111001;
		14'b11111100111011:	sigmoid = 21'b011001111010110010100;
		14'b11111100111100:	sigmoid = 21'b011001111100101101111;
		14'b11111100111101:	sigmoid = 21'b011001111110101001011;
		14'b11111100111110:	sigmoid = 21'b011010000000100100111;
		14'b11111100111111:	sigmoid = 21'b011010000010100000011;
		14'b11111101000000:	sigmoid = 21'b011010000100011100000;
		14'b11111101000001:	sigmoid = 21'b011010000110010111101;
		14'b11111101000010:	sigmoid = 21'b011010001000010011010;
		14'b11111101000011:	sigmoid = 21'b011010001010001111000;
		14'b11111101000100:	sigmoid = 21'b011010001100001010110;
		14'b11111101000101:	sigmoid = 21'b011010001110000110100;
		14'b11111101000110:	sigmoid = 21'b011010010000000010011;
		14'b11111101000111:	sigmoid = 21'b011010010001111110010;
		14'b11111101001000:	sigmoid = 21'b011010010011111010001;
		14'b11111101001001:	sigmoid = 21'b011010010101110110001;
		14'b11111101001010:	sigmoid = 21'b011010010111110010001;
		14'b11111101001011:	sigmoid = 21'b011010011001101110010;
		14'b11111101001100:	sigmoid = 21'b011010011011101010011;
		14'b11111101001101:	sigmoid = 21'b011010011101100110100;
		14'b11111101001110:	sigmoid = 21'b011010011111100010101;
		14'b11111101001111:	sigmoid = 21'b011010100001011110111;
		14'b11111101010000:	sigmoid = 21'b011010100011011011001;
		14'b11111101010001:	sigmoid = 21'b011010100101010111100;
		14'b11111101010010:	sigmoid = 21'b011010100111010011111;
		14'b11111101010011:	sigmoid = 21'b011010101001010000010;
		14'b11111101010100:	sigmoid = 21'b011010101011001100101;
		14'b11111101010101:	sigmoid = 21'b011010101101001001001;
		14'b11111101010110:	sigmoid = 21'b011010101111000101101;
		14'b11111101010111:	sigmoid = 21'b011010110001000010010;
		14'b11111101011000:	sigmoid = 21'b011010110010111110111;
		14'b11111101011001:	sigmoid = 21'b011010110100111011100;
		14'b11111101011010:	sigmoid = 21'b011010110110111000001;
		14'b11111101011011:	sigmoid = 21'b011010111000110100111;
		14'b11111101011100:	sigmoid = 21'b011010111010110001101;
		14'b11111101011101:	sigmoid = 21'b011010111100101110011;
		14'b11111101011110:	sigmoid = 21'b011010111110101011010;
		14'b11111101011111:	sigmoid = 21'b011011000000101000001;
		14'b11111101100000:	sigmoid = 21'b011011000010100101000;
		14'b11111101100001:	sigmoid = 21'b011011000100100001111;
		14'b11111101100010:	sigmoid = 21'b011011000110011110111;
		14'b11111101100011:	sigmoid = 21'b011011001000011011111;
		14'b11111101100100:	sigmoid = 21'b011011001010011001000;
		14'b11111101100101:	sigmoid = 21'b011011001100010110001;
		14'b11111101100110:	sigmoid = 21'b011011001110010011010;
		14'b11111101100111:	sigmoid = 21'b011011010000010000011;
		14'b11111101101000:	sigmoid = 21'b011011010010001101101;
		14'b11111101101001:	sigmoid = 21'b011011010100001010111;
		14'b11111101101010:	sigmoid = 21'b011011010110001000001;
		14'b11111101101011:	sigmoid = 21'b011011011000000101011;
		14'b11111101101100:	sigmoid = 21'b011011011010000010110;
		14'b11111101101101:	sigmoid = 21'b011011011100000000001;
		14'b11111101101110:	sigmoid = 21'b011011011101111101100;
		14'b11111101101111:	sigmoid = 21'b011011011111111011000;
		14'b11111101110000:	sigmoid = 21'b011011100001111000100;
		14'b11111101110001:	sigmoid = 21'b011011100011110110000;
		14'b11111101110010:	sigmoid = 21'b011011100101110011100;
		14'b11111101110011:	sigmoid = 21'b011011100111110001001;
		14'b11111101110100:	sigmoid = 21'b011011101001101110110;
		14'b11111101110101:	sigmoid = 21'b011011101011101100011;
		14'b11111101110110:	sigmoid = 21'b011011101101101010001;
		14'b11111101110111:	sigmoid = 21'b011011101111100111111;
		14'b11111101111000:	sigmoid = 21'b011011110001100101101;
		14'b11111101111001:	sigmoid = 21'b011011110011100011011;
		14'b11111101111010:	sigmoid = 21'b011011110101100001001;
		14'b11111101111011:	sigmoid = 21'b011011110111011111000;
		14'b11111101111100:	sigmoid = 21'b011011111001011100111;
		14'b11111101111101:	sigmoid = 21'b011011111011011010111;
		14'b11111101111110:	sigmoid = 21'b011011111101011000110;
		14'b11111101111111:	sigmoid = 21'b011011111111010110110;
		14'b11111110000000:	sigmoid = 21'b011100000001010100110;
		14'b11111110000001:	sigmoid = 21'b011100000011010010110;
		14'b11111110000010:	sigmoid = 21'b011100000101010000111;
		14'b11111110000011:	sigmoid = 21'b011100000111001111000;
		14'b11111110000100:	sigmoid = 21'b011100001001001101001;
		14'b11111110000101:	sigmoid = 21'b011100001011001011010;
		14'b11111110000110:	sigmoid = 21'b011100001101001001011;
		14'b11111110000111:	sigmoid = 21'b011100001111000111101;
		14'b11111110001000:	sigmoid = 21'b011100010001000101111;
		14'b11111110001001:	sigmoid = 21'b011100010011000100001;
		14'b11111110001010:	sigmoid = 21'b011100010101000010100;
		14'b11111110001011:	sigmoid = 21'b011100010111000000110;
		14'b11111110001100:	sigmoid = 21'b011100011000111111001;
		14'b11111110001101:	sigmoid = 21'b011100011010111101100;
		14'b11111110001110:	sigmoid = 21'b011100011100111011111;
		14'b11111110001111:	sigmoid = 21'b011100011110111010011;
		14'b11111110010000:	sigmoid = 21'b011100100000111000111;
		14'b11111110010001:	sigmoid = 21'b011100100010110111011;
		14'b11111110010010:	sigmoid = 21'b011100100100110101111;
		14'b11111110010011:	sigmoid = 21'b011100100110110100011;
		14'b11111110010100:	sigmoid = 21'b011100101000110011000;
		14'b11111110010101:	sigmoid = 21'b011100101010110001101;
		14'b11111110010110:	sigmoid = 21'b011100101100110000010;
		14'b11111110010111:	sigmoid = 21'b011100101110101110111;
		14'b11111110011000:	sigmoid = 21'b011100110000101101100;
		14'b11111110011001:	sigmoid = 21'b011100110010101100010;
		14'b11111110011010:	sigmoid = 21'b011100110100101011000;
		14'b11111110011011:	sigmoid = 21'b011100110110101001110;
		14'b11111110011100:	sigmoid = 21'b011100111000101000100;
		14'b11111110011101:	sigmoid = 21'b011100111010100111010;
		14'b11111110011110:	sigmoid = 21'b011100111100100110001;
		14'b11111110011111:	sigmoid = 21'b011100111110100101000;
		14'b11111110100000:	sigmoid = 21'b011101000000100011110;
		14'b11111110100001:	sigmoid = 21'b011101000010100010110;
		14'b11111110100010:	sigmoid = 21'b011101000100100001101;
		14'b11111110100011:	sigmoid = 21'b011101000110100000100;
		14'b11111110100100:	sigmoid = 21'b011101001000011111100;
		14'b11111110100101:	sigmoid = 21'b011101001010011110100;
		14'b11111110100110:	sigmoid = 21'b011101001100011101100;
		14'b11111110100111:	sigmoid = 21'b011101001110011100100;
		14'b11111110101000:	sigmoid = 21'b011101010000011011101;
		14'b11111110101001:	sigmoid = 21'b011101010010011010101;
		14'b11111110101010:	sigmoid = 21'b011101010100011001110;
		14'b11111110101011:	sigmoid = 21'b011101010110011000111;
		14'b11111110101100:	sigmoid = 21'b011101011000011000000;
		14'b11111110101101:	sigmoid = 21'b011101011010010111001;
		14'b11111110101110:	sigmoid = 21'b011101011100010110011;
		14'b11111110101111:	sigmoid = 21'b011101011110010101100;
		14'b11111110110000:	sigmoid = 21'b011101100000010100110;
		14'b11111110110001:	sigmoid = 21'b011101100010010100000;
		14'b11111110110010:	sigmoid = 21'b011101100100010011010;
		14'b11111110110011:	sigmoid = 21'b011101100110010010100;
		14'b11111110110100:	sigmoid = 21'b011101101000010001110;
		14'b11111110110101:	sigmoid = 21'b011101101010010001001;
		14'b11111110110110:	sigmoid = 21'b011101101100010000011;
		14'b11111110110111:	sigmoid = 21'b011101101110001111110;
		14'b11111110111000:	sigmoid = 21'b011101110000001111001;
		14'b11111110111001:	sigmoid = 21'b011101110010001110100;
		14'b11111110111010:	sigmoid = 21'b011101110100001101111;
		14'b11111110111011:	sigmoid = 21'b011101110110001101010;
		14'b11111110111100:	sigmoid = 21'b011101111000001100110;
		14'b11111110111101:	sigmoid = 21'b011101111010001100001;
		14'b11111110111110:	sigmoid = 21'b011101111100001011101;
		14'b11111110111111:	sigmoid = 21'b011101111110001011001;
		14'b11111111000000:	sigmoid = 21'b011110000000001010101;
		14'b11111111000001:	sigmoid = 21'b011110000010001010001;
		14'b11111111000010:	sigmoid = 21'b011110000100001001101;
		14'b11111111000011:	sigmoid = 21'b011110000110001001001;
		14'b11111111000100:	sigmoid = 21'b011110001000001000110;
		14'b11111111000101:	sigmoid = 21'b011110001010001000010;
		14'b11111111000110:	sigmoid = 21'b011110001100000111111;
		14'b11111111000111:	sigmoid = 21'b011110001110000111100;
		14'b11111111001000:	sigmoid = 21'b011110010000000111001;
		14'b11111111001001:	sigmoid = 21'b011110010010000110110;
		14'b11111111001010:	sigmoid = 21'b011110010100000110011;
		14'b11111111001011:	sigmoid = 21'b011110010110000110000;
		14'b11111111001100:	sigmoid = 21'b011110011000000101101;
		14'b11111111001101:	sigmoid = 21'b011110011010000101011;
		14'b11111111001110:	sigmoid = 21'b011110011100000101000;
		14'b11111111001111:	sigmoid = 21'b011110011110000100110;
		14'b11111111010000:	sigmoid = 21'b011110100000000100011;
		14'b11111111010001:	sigmoid = 21'b011110100010000100001;
		14'b11111111010010:	sigmoid = 21'b011110100100000011111;
		14'b11111111010011:	sigmoid = 21'b011110100110000011101;
		14'b11111111010100:	sigmoid = 21'b011110101000000011011;
		14'b11111111010101:	sigmoid = 21'b011110101010000011001;
		14'b11111111010110:	sigmoid = 21'b011110101100000011000;
		14'b11111111010111:	sigmoid = 21'b011110101110000010110;
		14'b11111111011000:	sigmoid = 21'b011110110000000010100;
		14'b11111111011001:	sigmoid = 21'b011110110010000010011;
		14'b11111111011010:	sigmoid = 21'b011110110100000010001;
		14'b11111111011011:	sigmoid = 21'b011110110110000010000;
		14'b11111111011100:	sigmoid = 21'b011110111000000001111;
		14'b11111111011101:	sigmoid = 21'b011110111010000001101;
		14'b11111111011110:	sigmoid = 21'b011110111100000001100;
		14'b11111111011111:	sigmoid = 21'b011110111110000001011;
		14'b11111111100000:	sigmoid = 21'b011111000000000001010;
		14'b11111111100001:	sigmoid = 21'b011111000010000001001;
		14'b11111111100010:	sigmoid = 21'b011111000100000001000;
		14'b11111111100011:	sigmoid = 21'b011111000110000000111;
		14'b11111111100100:	sigmoid = 21'b011111001000000000111;
		14'b11111111100101:	sigmoid = 21'b011111001010000000110;
		14'b11111111100110:	sigmoid = 21'b011111001100000000101;
		14'b11111111100111:	sigmoid = 21'b011111001110000000101;
		14'b11111111101000:	sigmoid = 21'b011111010000000000100;
		14'b11111111101001:	sigmoid = 21'b011111010010000000011;
		14'b11111111101010:	sigmoid = 21'b011111010100000000011;
		14'b11111111101011:	sigmoid = 21'b011111010110000000011;
		14'b11111111101100:	sigmoid = 21'b011111011000000000010;
		14'b11111111101101:	sigmoid = 21'b011111011010000000010;
		14'b11111111101110:	sigmoid = 21'b011111011100000000001;
		14'b11111111101111:	sigmoid = 21'b011111011110000000001;
		14'b11111111110000:	sigmoid = 21'b011111100000000000001;
		14'b11111111110001:	sigmoid = 21'b011111100010000000001;
		14'b11111111110010:	sigmoid = 21'b011111100100000000000;
		14'b11111111110011:	sigmoid = 21'b011111100110000000000;
		14'b11111111110100:	sigmoid = 21'b011111101000000000000;
		14'b11111111110101:	sigmoid = 21'b011111101010000000000;
		14'b11111111110110:	sigmoid = 21'b011111101100000000000;
		14'b11111111110111:	sigmoid = 21'b011111101110000000000;
		14'b11111111111000:	sigmoid = 21'b011111110000000000000;
		14'b11111111111001:	sigmoid = 21'b011111110010000000000;
		14'b11111111111010:	sigmoid = 21'b011111110100000000000;
		14'b11111111111011:	sigmoid = 21'b011111110110000000000;
		14'b11111111111100:	sigmoid = 21'b011111111000000000000;
		14'b11111111111101:	sigmoid = 21'b011111111010000000000;
		14'b11111111111110:	sigmoid = 21'b011111111100000000000;
		14'b11111111111111:	sigmoid = 21'b011111111110000000000;
		14'b00000000000000:	sigmoid = 21'b100000000000000000000;
		14'b00000000000001:	sigmoid = 21'b100000000001111111111;
		14'b00000000000010:	sigmoid = 21'b100000000011111111111;
		14'b00000000000011:	sigmoid = 21'b100000000101111111111;
		14'b00000000000100:	sigmoid = 21'b100000000111111111111;
		14'b00000000000101:	sigmoid = 21'b100000001001111111111;
		14'b00000000000110:	sigmoid = 21'b100000001011111111111;
		14'b00000000000111:	sigmoid = 21'b100000001101111111111;
		14'b00000000001000:	sigmoid = 21'b100000001111111111111;
		14'b00000000001001:	sigmoid = 21'b100000010001111111111;
		14'b00000000001010:	sigmoid = 21'b100000010011111111111;
		14'b00000000001011:	sigmoid = 21'b100000010101111111111;
		14'b00000000001100:	sigmoid = 21'b100000010111111111111;
		14'b00000000001101:	sigmoid = 21'b100000011001111111111;
		14'b00000000001110:	sigmoid = 21'b100000011011111111111;
		14'b00000000001111:	sigmoid = 21'b100000011101111111110;
		14'b00000000010000:	sigmoid = 21'b100000011111111111110;
		14'b00000000010001:	sigmoid = 21'b100000100001111111110;
		14'b00000000010010:	sigmoid = 21'b100000100011111111110;
		14'b00000000010011:	sigmoid = 21'b100000100101111111101;
		14'b00000000010100:	sigmoid = 21'b100000100111111111101;
		14'b00000000010101:	sigmoid = 21'b100000101001111111100;
		14'b00000000010110:	sigmoid = 21'b100000101011111111100;
		14'b00000000010111:	sigmoid = 21'b100000101101111111100;
		14'b00000000011000:	sigmoid = 21'b100000101111111111011;
		14'b00000000011001:	sigmoid = 21'b100000110001111111010;
		14'b00000000011010:	sigmoid = 21'b100000110011111111010;
		14'b00000000011011:	sigmoid = 21'b100000110101111111001;
		14'b00000000011100:	sigmoid = 21'b100000110111111111000;
		14'b00000000011101:	sigmoid = 21'b100000111001111111000;
		14'b00000000011110:	sigmoid = 21'b100000111011111110111;
		14'b00000000011111:	sigmoid = 21'b100000111101111110110;
		14'b00000000100000:	sigmoid = 21'b100000111111111110101;
		14'b00000000100001:	sigmoid = 21'b100001000001111110100;
		14'b00000000100010:	sigmoid = 21'b100001000011111110011;
		14'b00000000100011:	sigmoid = 21'b100001000101111110010;
		14'b00000000100100:	sigmoid = 21'b100001000111111110000;
		14'b00000000100101:	sigmoid = 21'b100001001001111101111;
		14'b00000000100110:	sigmoid = 21'b100001001011111101110;
		14'b00000000100111:	sigmoid = 21'b100001001101111101100;
		14'b00000000101000:	sigmoid = 21'b100001001111111101011;
		14'b00000000101001:	sigmoid = 21'b100001010001111101001;
		14'b00000000101010:	sigmoid = 21'b100001010011111100111;
		14'b00000000101011:	sigmoid = 21'b100001010101111100110;
		14'b00000000101100:	sigmoid = 21'b100001010111111100100;
		14'b00000000101101:	sigmoid = 21'b100001011001111100010;
		14'b00000000101110:	sigmoid = 21'b100001011011111100000;
		14'b00000000101111:	sigmoid = 21'b100001011101111011110;
		14'b00000000110000:	sigmoid = 21'b100001011111111011100;
		14'b00000000110001:	sigmoid = 21'b100001100001111011001;
		14'b00000000110010:	sigmoid = 21'b100001100011111010111;
		14'b00000000110011:	sigmoid = 21'b100001100101111010100;
		14'b00000000110100:	sigmoid = 21'b100001100111111010010;
		14'b00000000110101:	sigmoid = 21'b100001101001111001111;
		14'b00000000110110:	sigmoid = 21'b100001101011111001100;
		14'b00000000110111:	sigmoid = 21'b100001101101111001001;
		14'b00000000111000:	sigmoid = 21'b100001101111111000110;
		14'b00000000111001:	sigmoid = 21'b100001110001111000011;
		14'b00000000111010:	sigmoid = 21'b100001110011111000000;
		14'b00000000111011:	sigmoid = 21'b100001110101110111101;
		14'b00000000111100:	sigmoid = 21'b100001110111110111001;
		14'b00000000111101:	sigmoid = 21'b100001111001110110110;
		14'b00000000111110:	sigmoid = 21'b100001111011110110010;
		14'b00000000111111:	sigmoid = 21'b100001111101110101110;
		14'b00000001000000:	sigmoid = 21'b100001111111110101010;
		14'b00000001000001:	sigmoid = 21'b100010000001110100110;
		14'b00000001000010:	sigmoid = 21'b100010000011110100010;
		14'b00000001000011:	sigmoid = 21'b100010000101110011110;
		14'b00000001000100:	sigmoid = 21'b100010000111110011001;
		14'b00000001000101:	sigmoid = 21'b100010001001110010101;
		14'b00000001000110:	sigmoid = 21'b100010001011110010000;
		14'b00000001000111:	sigmoid = 21'b100010001101110001011;
		14'b00000001001000:	sigmoid = 21'b100010001111110000110;
		14'b00000001001001:	sigmoid = 21'b100010010001110000001;
		14'b00000001001010:	sigmoid = 21'b100010010011101111100;
		14'b00000001001011:	sigmoid = 21'b100010010101101110110;
		14'b00000001001100:	sigmoid = 21'b100010010111101110001;
		14'b00000001001101:	sigmoid = 21'b100010011001101101011;
		14'b00000001001110:	sigmoid = 21'b100010011011101100101;
		14'b00000001001111:	sigmoid = 21'b100010011101101011111;
		14'b00000001010000:	sigmoid = 21'b100010011111101011001;
		14'b00000001010001:	sigmoid = 21'b100010100001101010011;
		14'b00000001010010:	sigmoid = 21'b100010100011101001100;
		14'b00000001010011:	sigmoid = 21'b100010100101101000110;
		14'b00000001010100:	sigmoid = 21'b100010100111100111111;
		14'b00000001010101:	sigmoid = 21'b100010101001100111000;
		14'b00000001010110:	sigmoid = 21'b100010101011100110001;
		14'b00000001010111:	sigmoid = 21'b100010101101100101010;
		14'b00000001011000:	sigmoid = 21'b100010101111100100010;
		14'b00000001011001:	sigmoid = 21'b100010110001100011011;
		14'b00000001011010:	sigmoid = 21'b100010110011100010011;
		14'b00000001011011:	sigmoid = 21'b100010110101100001011;
		14'b00000001011100:	sigmoid = 21'b100010110111100000011;
		14'b00000001011101:	sigmoid = 21'b100010111001011111011;
		14'b00000001011110:	sigmoid = 21'b100010111011011110010;
		14'b00000001011111:	sigmoid = 21'b100010111101011101001;
		14'b00000001100000:	sigmoid = 21'b100010111111011100001;
		14'b00000001100001:	sigmoid = 21'b100011000001011010111;
		14'b00000001100010:	sigmoid = 21'b100011000011011001110;
		14'b00000001100011:	sigmoid = 21'b100011000101011000101;
		14'b00000001100100:	sigmoid = 21'b100011000111010111011;
		14'b00000001100101:	sigmoid = 21'b100011001001010110001;
		14'b00000001100110:	sigmoid = 21'b100011001011010100111;
		14'b00000001100111:	sigmoid = 21'b100011001101010011101;
		14'b00000001101000:	sigmoid = 21'b100011001111010010011;
		14'b00000001101001:	sigmoid = 21'b100011010001010001000;
		14'b00000001101010:	sigmoid = 21'b100011010011001111101;
		14'b00000001101011:	sigmoid = 21'b100011010101001110010;
		14'b00000001101100:	sigmoid = 21'b100011010111001100111;
		14'b00000001101101:	sigmoid = 21'b100011011001001011100;
		14'b00000001101110:	sigmoid = 21'b100011011011001010000;
		14'b00000001101111:	sigmoid = 21'b100011011101001000100;
		14'b00000001110000:	sigmoid = 21'b100011011111000111000;
		14'b00000001110001:	sigmoid = 21'b100011100001000101100;
		14'b00000001110010:	sigmoid = 21'b100011100011000100000;
		14'b00000001110011:	sigmoid = 21'b100011100101000010011;
		14'b00000001110100:	sigmoid = 21'b100011100111000000110;
		14'b00000001110101:	sigmoid = 21'b100011101000111111001;
		14'b00000001110110:	sigmoid = 21'b100011101010111101011;
		14'b00000001110111:	sigmoid = 21'b100011101100111011110;
		14'b00000001111000:	sigmoid = 21'b100011101110111010000;
		14'b00000001111001:	sigmoid = 21'b100011110000111000010;
		14'b00000001111010:	sigmoid = 21'b100011110010110110100;
		14'b00000001111011:	sigmoid = 21'b100011110100110100101;
		14'b00000001111100:	sigmoid = 21'b100011110110110010110;
		14'b00000001111101:	sigmoid = 21'b100011111000110000111;
		14'b00000001111110:	sigmoid = 21'b100011111010101111000;
		14'b00000001111111:	sigmoid = 21'b100011111100101101001;
		14'b00000010000000:	sigmoid = 21'b100011111110101011001;
		14'b00000010000001:	sigmoid = 21'b100100000000101001001;
		14'b00000010000010:	sigmoid = 21'b100100000010100111001;
		14'b00000010000011:	sigmoid = 21'b100100000100100101000;
		14'b00000010000100:	sigmoid = 21'b100100000110100011000;
		14'b00000010000101:	sigmoid = 21'b100100001000100000111;
		14'b00000010000110:	sigmoid = 21'b100100001010011110110;
		14'b00000010000111:	sigmoid = 21'b100100001100011100100;
		14'b00000010001000:	sigmoid = 21'b100100001110011010010;
		14'b00000010001001:	sigmoid = 21'b100100010000011000000;
		14'b00000010001010:	sigmoid = 21'b100100010010010101110;
		14'b00000010001011:	sigmoid = 21'b100100010100010011100;
		14'b00000010001100:	sigmoid = 21'b100100010110010001001;
		14'b00000010001101:	sigmoid = 21'b100100011000001110110;
		14'b00000010001110:	sigmoid = 21'b100100011010001100011;
		14'b00000010001111:	sigmoid = 21'b100100011100001001111;
		14'b00000010010000:	sigmoid = 21'b100100011110000111011;
		14'b00000010010001:	sigmoid = 21'b100100100000000100111;
		14'b00000010010010:	sigmoid = 21'b100100100010000010011;
		14'b00000010010011:	sigmoid = 21'b100100100011111111110;
		14'b00000010010100:	sigmoid = 21'b100100100101111101001;
		14'b00000010010101:	sigmoid = 21'b100100100111111010100;
		14'b00000010010110:	sigmoid = 21'b100100101001110111110;
		14'b00000010010111:	sigmoid = 21'b100100101011110101000;
		14'b00000010011000:	sigmoid = 21'b100100101101110010010;
		14'b00000010011001:	sigmoid = 21'b100100101111101111100;
		14'b00000010011010:	sigmoid = 21'b100100110001101100101;
		14'b00000010011011:	sigmoid = 21'b100100110011101001110;
		14'b00000010011100:	sigmoid = 21'b100100110101100110111;
		14'b00000010011101:	sigmoid = 21'b100100110111100100000;
		14'b00000010011110:	sigmoid = 21'b100100111001100001000;
		14'b00000010011111:	sigmoid = 21'b100100111011011110000;
		14'b00000010100000:	sigmoid = 21'b100100111101011010111;
		14'b00000010100001:	sigmoid = 21'b100100111111010111110;
		14'b00000010100010:	sigmoid = 21'b100101000001010100101;
		14'b00000010100011:	sigmoid = 21'b100101000011010001100;
		14'b00000010100100:	sigmoid = 21'b100101000101001110010;
		14'b00000010100101:	sigmoid = 21'b100101000111001011000;
		14'b00000010100110:	sigmoid = 21'b100101001001000111110;
		14'b00000010100111:	sigmoid = 21'b100101001011000100011;
		14'b00000010101000:	sigmoid = 21'b100101001101000001000;
		14'b00000010101001:	sigmoid = 21'b100101001110111101101;
		14'b00000010101010:	sigmoid = 21'b100101010000111010010;
		14'b00000010101011:	sigmoid = 21'b100101010010110110110;
		14'b00000010101100:	sigmoid = 21'b100101010100110011010;
		14'b00000010101101:	sigmoid = 21'b100101010110101111101;
		14'b00000010101110:	sigmoid = 21'b100101011000101100000;
		14'b00000010101111:	sigmoid = 21'b100101011010101000011;
		14'b00000010110000:	sigmoid = 21'b100101011100100100110;
		14'b00000010110001:	sigmoid = 21'b100101011110100001000;
		14'b00000010110010:	sigmoid = 21'b100101100000011101010;
		14'b00000010110011:	sigmoid = 21'b100101100010011001011;
		14'b00000010110100:	sigmoid = 21'b100101100100010101100;
		14'b00000010110101:	sigmoid = 21'b100101100110010001101;
		14'b00000010110110:	sigmoid = 21'b100101101000001101110;
		14'b00000010110111:	sigmoid = 21'b100101101010001001110;
		14'b00000010111000:	sigmoid = 21'b100101101100000101110;
		14'b00000010111001:	sigmoid = 21'b100101101110000001101;
		14'b00000010111010:	sigmoid = 21'b100101101111111101100;
		14'b00000010111011:	sigmoid = 21'b100101110001111001011;
		14'b00000010111100:	sigmoid = 21'b100101110011110101001;
		14'b00000010111101:	sigmoid = 21'b100101110101110000111;
		14'b00000010111110:	sigmoid = 21'b100101110111101100101;
		14'b00000010111111:	sigmoid = 21'b100101111001101000010;
		14'b00000011000000:	sigmoid = 21'b100101111011100011111;
		14'b00000011000001:	sigmoid = 21'b100101111101011111100;
		14'b00000011000010:	sigmoid = 21'b100101111111011011000;
		14'b00000011000011:	sigmoid = 21'b100110000001010110100;
		14'b00000011000100:	sigmoid = 21'b100110000011010010000;
		14'b00000011000101:	sigmoid = 21'b100110000101001101011;
		14'b00000011000110:	sigmoid = 21'b100110000111001000110;
		14'b00000011000111:	sigmoid = 21'b100110001001000100000;
		14'b00000011001000:	sigmoid = 21'b100110001010111111010;
		14'b00000011001001:	sigmoid = 21'b100110001100111010100;
		14'b00000011001010:	sigmoid = 21'b100110001110110101110;
		14'b00000011001011:	sigmoid = 21'b100110010000110000111;
		14'b00000011001100:	sigmoid = 21'b100110010010101011111;
		14'b00000011001101:	sigmoid = 21'b100110010100100110111;
		14'b00000011001110:	sigmoid = 21'b100110010110100001111;
		14'b00000011001111:	sigmoid = 21'b100110011000011100111;
		14'b00000011010000:	sigmoid = 21'b100110011010010111110;
		14'b00000011010001:	sigmoid = 21'b100110011100010010100;
		14'b00000011010010:	sigmoid = 21'b100110011110001101011;
		14'b00000011010011:	sigmoid = 21'b100110100000001000001;
		14'b00000011010100:	sigmoid = 21'b100110100010000010110;
		14'b00000011010101:	sigmoid = 21'b100110100011111101011;
		14'b00000011010110:	sigmoid = 21'b100110100101111000000;
		14'b00000011010111:	sigmoid = 21'b100110100111110010100;
		14'b00000011011000:	sigmoid = 21'b100110101001101101000;
		14'b00000011011001:	sigmoid = 21'b100110101011100111100;
		14'b00000011011010:	sigmoid = 21'b100110101101100001111;
		14'b00000011011011:	sigmoid = 21'b100110101111011100010;
		14'b00000011011100:	sigmoid = 21'b100110110001010110100;
		14'b00000011011101:	sigmoid = 21'b100110110011010000110;
		14'b00000011011110:	sigmoid = 21'b100110110101001011000;
		14'b00000011011111:	sigmoid = 21'b100110110111000101001;
		14'b00000011100000:	sigmoid = 21'b100110111000111111010;
		14'b00000011100001:	sigmoid = 21'b100110111010111001010;
		14'b00000011100010:	sigmoid = 21'b100110111100110011010;
		14'b00000011100011:	sigmoid = 21'b100110111110101101001;
		14'b00000011100100:	sigmoid = 21'b100111000000100111000;
		14'b00000011100101:	sigmoid = 21'b100111000010100000111;
		14'b00000011100110:	sigmoid = 21'b100111000100011010101;
		14'b00000011100111:	sigmoid = 21'b100111000110010100011;
		14'b00000011101000:	sigmoid = 21'b100111001000001110000;
		14'b00000011101001:	sigmoid = 21'b100111001010000111101;
		14'b00000011101010:	sigmoid = 21'b100111001100000001010;
		14'b00000011101011:	sigmoid = 21'b100111001101111010110;
		14'b00000011101100:	sigmoid = 21'b100111001111110100010;
		14'b00000011101101:	sigmoid = 21'b100111010001101101101;
		14'b00000011101110:	sigmoid = 21'b100111010011100111000;
		14'b00000011101111:	sigmoid = 21'b100111010101100000010;
		14'b00000011110000:	sigmoid = 21'b100111010111011001100;
		14'b00000011110001:	sigmoid = 21'b100111011001010010110;
		14'b00000011110010:	sigmoid = 21'b100111011011001011111;
		14'b00000011110011:	sigmoid = 21'b100111011101000101000;
		14'b00000011110100:	sigmoid = 21'b100111011110111110000;
		14'b00000011110101:	sigmoid = 21'b100111100000110110111;
		14'b00000011110110:	sigmoid = 21'b100111100010101111111;
		14'b00000011110111:	sigmoid = 21'b100111100100101000110;
		14'b00000011111000:	sigmoid = 21'b100111100110100001100;
		14'b00000011111001:	sigmoid = 21'b100111101000011010010;
		14'b00000011111010:	sigmoid = 21'b100111101010010011000;
		14'b00000011111011:	sigmoid = 21'b100111101100001011101;
		14'b00000011111100:	sigmoid = 21'b100111101110000100001;
		14'b00000011111101:	sigmoid = 21'b100111101111111100110;
		14'b00000011111110:	sigmoid = 21'b100111110001110101001;
		14'b00000011111111:	sigmoid = 21'b100111110011101101101;
		14'b00000100000000:	sigmoid = 21'b100111110101100101111;
		14'b00000100000001:	sigmoid = 21'b100111110111011110010;
		14'b00000100000010:	sigmoid = 21'b100111111001010110100;
		14'b00000100000011:	sigmoid = 21'b100111111011001110101;
		14'b00000100000100:	sigmoid = 21'b100111111101000110110;
		14'b00000100000101:	sigmoid = 21'b100111111110111110110;
		14'b00000100000110:	sigmoid = 21'b101000000000110110110;
		14'b00000100000111:	sigmoid = 21'b101000000010101110110;
		14'b00000100001000:	sigmoid = 21'b101000000100100110101;
		14'b00000100001001:	sigmoid = 21'b101000000110011110100;
		14'b00000100001010:	sigmoid = 21'b101000001000010110010;
		14'b00000100001011:	sigmoid = 21'b101000001010001101111;
		14'b00000100001100:	sigmoid = 21'b101000001100000101101;
		14'b00000100001101:	sigmoid = 21'b101000001101111101001;
		14'b00000100001110:	sigmoid = 21'b101000001111110100110;
		14'b00000100001111:	sigmoid = 21'b101000010001101100001;
		14'b00000100010000:	sigmoid = 21'b101000010011100011101;
		14'b00000100010001:	sigmoid = 21'b101000010101011010111;
		14'b00000100010010:	sigmoid = 21'b101000010111010010010;
		14'b00000100010011:	sigmoid = 21'b101000011001001001011;
		14'b00000100010100:	sigmoid = 21'b101000011011000000101;
		14'b00000100010101:	sigmoid = 21'b101000011100110111110;
		14'b00000100010110:	sigmoid = 21'b101000011110101110110;
		14'b00000100010111:	sigmoid = 21'b101000100000100101110;
		14'b00000100011000:	sigmoid = 21'b101000100010011100101;
		14'b00000100011001:	sigmoid = 21'b101000100100010011100;
		14'b00000100011010:	sigmoid = 21'b101000100110001010010;
		14'b00000100011011:	sigmoid = 21'b101000101000000001000;
		14'b00000100011100:	sigmoid = 21'b101000101001110111110;
		14'b00000100011101:	sigmoid = 21'b101000101011101110010;
		14'b00000100011110:	sigmoid = 21'b101000101101100100111;
		14'b00000100011111:	sigmoid = 21'b101000101111011011011;
		14'b00000100100000:	sigmoid = 21'b101000110001010001110;
		14'b00000100100001:	sigmoid = 21'b101000110011001000001;
		14'b00000100100010:	sigmoid = 21'b101000110100111110011;
		14'b00000100100011:	sigmoid = 21'b101000110110110100101;
		14'b00000100100100:	sigmoid = 21'b101000111000101010110;
		14'b00000100100101:	sigmoid = 21'b101000111010100000111;
		14'b00000100100110:	sigmoid = 21'b101000111100010110111;
		14'b00000100100111:	sigmoid = 21'b101000111110001100111;
		14'b00000100101000:	sigmoid = 21'b101001000000000010110;
		14'b00000100101001:	sigmoid = 21'b101001000001111000101;
		14'b00000100101010:	sigmoid = 21'b101001000011101110011;
		14'b00000100101011:	sigmoid = 21'b101001000101100100001;
		14'b00000100101100:	sigmoid = 21'b101001000111011001110;
		14'b00000100101101:	sigmoid = 21'b101001001001001111011;
		14'b00000100101110:	sigmoid = 21'b101001001011000100111;
		14'b00000100101111:	sigmoid = 21'b101001001100111010010;
		14'b00000100110000:	sigmoid = 21'b101001001110101111101;
		14'b00000100110001:	sigmoid = 21'b101001010000100101000;
		14'b00000100110010:	sigmoid = 21'b101001010010011010010;
		14'b00000100110011:	sigmoid = 21'b101001010100001111011;
		14'b00000100110100:	sigmoid = 21'b101001010110000100100;
		14'b00000100110101:	sigmoid = 21'b101001010111111001101;
		14'b00000100110110:	sigmoid = 21'b101001011001101110101;
		14'b00000100110111:	sigmoid = 21'b101001011011100011100;
		14'b00000100111000:	sigmoid = 21'b101001011101011000011;
		14'b00000100111001:	sigmoid = 21'b101001011111001101001;
		14'b00000100111010:	sigmoid = 21'b101001100001000001111;
		14'b00000100111011:	sigmoid = 21'b101001100010110110100;
		14'b00000100111100:	sigmoid = 21'b101001100100101011001;
		14'b00000100111101:	sigmoid = 21'b101001100110011111101;
		14'b00000100111110:	sigmoid = 21'b101001101000010100000;
		14'b00000100111111:	sigmoid = 21'b101001101010001000011;
		14'b00000101000000:	sigmoid = 21'b101001101011111100110;
		14'b00000101000001:	sigmoid = 21'b101001101101110001000;
		14'b00000101000010:	sigmoid = 21'b101001101111100101001;
		14'b00000101000011:	sigmoid = 21'b101001110001011001010;
		14'b00000101000100:	sigmoid = 21'b101001110011001101010;
		14'b00000101000101:	sigmoid = 21'b101001110101000001010;
		14'b00000101000110:	sigmoid = 21'b101001110110110101001;
		14'b00000101000111:	sigmoid = 21'b101001111000101000111;
		14'b00000101001000:	sigmoid = 21'b101001111010011100101;
		14'b00000101001001:	sigmoid = 21'b101001111100010000011;
		14'b00000101001010:	sigmoid = 21'b101001111110000100000;
		14'b00000101001011:	sigmoid = 21'b101001111111110111100;
		14'b00000101001100:	sigmoid = 21'b101010000001101011000;
		14'b00000101001101:	sigmoid = 21'b101010000011011110011;
		14'b00000101001110:	sigmoid = 21'b101010000101010001110;
		14'b00000101001111:	sigmoid = 21'b101010000111000101000;
		14'b00000101010000:	sigmoid = 21'b101010001000111000001;
		14'b00000101010001:	sigmoid = 21'b101010001010101011010;
		14'b00000101010010:	sigmoid = 21'b101010001100011110010;
		14'b00000101010011:	sigmoid = 21'b101010001110010001010;
		14'b00000101010100:	sigmoid = 21'b101010010000000100001;
		14'b00000101010101:	sigmoid = 21'b101010010001110111000;
		14'b00000101010110:	sigmoid = 21'b101010010011101001110;
		14'b00000101010111:	sigmoid = 21'b101010010101011100011;
		14'b00000101011000:	sigmoid = 21'b101010010111001111000;
		14'b00000101011001:	sigmoid = 21'b101010011001000001101;
		14'b00000101011010:	sigmoid = 21'b101010011010110100000;
		14'b00000101011011:	sigmoid = 21'b101010011100100110100;
		14'b00000101011100:	sigmoid = 21'b101010011110011000110;
		14'b00000101011101:	sigmoid = 21'b101010100000001011000;
		14'b00000101011110:	sigmoid = 21'b101010100001111101010;
		14'b00000101011111:	sigmoid = 21'b101010100011101111010;
		14'b00000101100000:	sigmoid = 21'b101010100101100001011;
		14'b00000101100001:	sigmoid = 21'b101010100111010011010;
		14'b00000101100010:	sigmoid = 21'b101010101001000101001;
		14'b00000101100011:	sigmoid = 21'b101010101010110111000;
		14'b00000101100100:	sigmoid = 21'b101010101100101000110;
		14'b00000101100101:	sigmoid = 21'b101010101110011010011;
		14'b00000101100110:	sigmoid = 21'b101010110000001100000;
		14'b00000101100111:	sigmoid = 21'b101010110001111101100;
		14'b00000101101000:	sigmoid = 21'b101010110011101110111;
		14'b00000101101001:	sigmoid = 21'b101010110101100000010;
		14'b00000101101010:	sigmoid = 21'b101010110111010001100;
		14'b00000101101011:	sigmoid = 21'b101010111001000010110;
		14'b00000101101100:	sigmoid = 21'b101010111010110011111;
		14'b00000101101101:	sigmoid = 21'b101010111100100100111;
		14'b00000101101110:	sigmoid = 21'b101010111110010101111;
		14'b00000101101111:	sigmoid = 21'b101011000000000110111;
		14'b00000101110000:	sigmoid = 21'b101011000001110111101;
		14'b00000101110001:	sigmoid = 21'b101011000011101000011;
		14'b00000101110010:	sigmoid = 21'b101011000101011001001;
		14'b00000101110011:	sigmoid = 21'b101011000111001001110;
		14'b00000101110100:	sigmoid = 21'b101011001000111010010;
		14'b00000101110101:	sigmoid = 21'b101011001010101010101;
		14'b00000101110110:	sigmoid = 21'b101011001100011011000;
		14'b00000101110111:	sigmoid = 21'b101011001110001011011;
		14'b00000101111000:	sigmoid = 21'b101011001111111011101;
		14'b00000101111001:	sigmoid = 21'b101011010001101011110;
		14'b00000101111010:	sigmoid = 21'b101011010011011011110;
		14'b00000101111011:	sigmoid = 21'b101011010101001011110;
		14'b00000101111100:	sigmoid = 21'b101011010110111011101;
		14'b00000101111101:	sigmoid = 21'b101011011000101011100;
		14'b00000101111110:	sigmoid = 21'b101011011010011011010;
		14'b00000101111111:	sigmoid = 21'b101011011100001011000;
		14'b00000110000000:	sigmoid = 21'b101011011101111010100;
		14'b00000110000001:	sigmoid = 21'b101011011111101010001;
		14'b00000110000010:	sigmoid = 21'b101011100001011001100;
		14'b00000110000011:	sigmoid = 21'b101011100011001000111;
		14'b00000110000100:	sigmoid = 21'b101011100100111000001;
		14'b00000110000101:	sigmoid = 21'b101011100110100111011;
		14'b00000110000110:	sigmoid = 21'b101011101000010110100;
		14'b00000110000111:	sigmoid = 21'b101011101010000101101;
		14'b00000110001000:	sigmoid = 21'b101011101011110100100;
		14'b00000110001001:	sigmoid = 21'b101011101101100011100;
		14'b00000110001010:	sigmoid = 21'b101011101111010010010;
		14'b00000110001011:	sigmoid = 21'b101011110001000001000;
		14'b00000110001100:	sigmoid = 21'b101011110010101111101;
		14'b00000110001101:	sigmoid = 21'b101011110100011110010;
		14'b00000110001110:	sigmoid = 21'b101011110110001100110;
		14'b00000110001111:	sigmoid = 21'b101011110111111011001;
		14'b00000110010000:	sigmoid = 21'b101011111001101001100;
		14'b00000110010001:	sigmoid = 21'b101011111011010111110;
		14'b00000110010010:	sigmoid = 21'b101011111101000101111;
		14'b00000110010011:	sigmoid = 21'b101011111110110100000;
		14'b00000110010100:	sigmoid = 21'b101100000000100010000;
		14'b00000110010101:	sigmoid = 21'b101100000010010000000;
		14'b00000110010110:	sigmoid = 21'b101100000011111101110;
		14'b00000110010111:	sigmoid = 21'b101100000101101011101;
		14'b00000110011000:	sigmoid = 21'b101100000111011001010;
		14'b00000110011001:	sigmoid = 21'b101100001001000110111;
		14'b00000110011010:	sigmoid = 21'b101100001010110100011;
		14'b00000110011011:	sigmoid = 21'b101100001100100001111;
		14'b00000110011100:	sigmoid = 21'b101100001110001111010;
		14'b00000110011101:	sigmoid = 21'b101100001111111100100;
		14'b00000110011110:	sigmoid = 21'b101100010001101001110;
		14'b00000110011111:	sigmoid = 21'b101100010011010110111;
		14'b00000110100000:	sigmoid = 21'b101100010101000011111;
		14'b00000110100001:	sigmoid = 21'b101100010110110000111;
		14'b00000110100010:	sigmoid = 21'b101100011000011101110;
		14'b00000110100011:	sigmoid = 21'b101100011010001010100;
		14'b00000110100100:	sigmoid = 21'b101100011011110111010;
		14'b00000110100101:	sigmoid = 21'b101100011101100011111;
		14'b00000110100110:	sigmoid = 21'b101100011111010000011;
		14'b00000110100111:	sigmoid = 21'b101100100000111100111;
		14'b00000110101000:	sigmoid = 21'b101100100010101001010;
		14'b00000110101001:	sigmoid = 21'b101100100100010101100;
		14'b00000110101010:	sigmoid = 21'b101100100110000001110;
		14'b00000110101011:	sigmoid = 21'b101100100111101101111;
		14'b00000110101100:	sigmoid = 21'b101100101001011001111;
		14'b00000110101101:	sigmoid = 21'b101100101011000101111;
		14'b00000110101110:	sigmoid = 21'b101100101100110001110;
		14'b00000110101111:	sigmoid = 21'b101100101110011101101;
		14'b00000110110000:	sigmoid = 21'b101100110000001001010;
		14'b00000110110001:	sigmoid = 21'b101100110001110100111;
		14'b00000110110010:	sigmoid = 21'b101100110011100000100;
		14'b00000110110011:	sigmoid = 21'b101100110101001011111;
		14'b00000110110100:	sigmoid = 21'b101100110110110111010;
		14'b00000110110101:	sigmoid = 21'b101100111000100010101;
		14'b00000110110110:	sigmoid = 21'b101100111010001101110;
		14'b00000110110111:	sigmoid = 21'b101100111011111000111;
		14'b00000110111000:	sigmoid = 21'b101100111101100100000;
		14'b00000110111001:	sigmoid = 21'b101100111111001110111;
		14'b00000110111010:	sigmoid = 21'b101101000000111001110;
		14'b00000110111011:	sigmoid = 21'b101101000010100100101;
		14'b00000110111100:	sigmoid = 21'b101101000100001111010;
		14'b00000110111101:	sigmoid = 21'b101101000101111001111;
		14'b00000110111110:	sigmoid = 21'b101101000111100100100;
		14'b00000110111111:	sigmoid = 21'b101101001001001110111;
		14'b00000111000000:	sigmoid = 21'b101101001010111001010;
		14'b00000111000001:	sigmoid = 21'b101101001100100011100;
		14'b00000111000010:	sigmoid = 21'b101101001110001101110;
		14'b00000111000011:	sigmoid = 21'b101101001111110111111;
		14'b00000111000100:	sigmoid = 21'b101101010001100001111;
		14'b00000111000101:	sigmoid = 21'b101101010011001011110;
		14'b00000111000110:	sigmoid = 21'b101101010100110101101;
		14'b00000111000111:	sigmoid = 21'b101101010110011111011;
		14'b00000111001000:	sigmoid = 21'b101101011000001001000;
		14'b00000111001001:	sigmoid = 21'b101101011001110010101;
		14'b00000111001010:	sigmoid = 21'b101101011011011100001;
		14'b00000111001011:	sigmoid = 21'b101101011101000101100;
		14'b00000111001100:	sigmoid = 21'b101101011110101110111;
		14'b00000111001101:	sigmoid = 21'b101101100000011000001;
		14'b00000111001110:	sigmoid = 21'b101101100010000001010;
		14'b00000111001111:	sigmoid = 21'b101101100011101010011;
		14'b00000111010000:	sigmoid = 21'b101101100101010011011;
		14'b00000111010001:	sigmoid = 21'b101101100110111100010;
		14'b00000111010010:	sigmoid = 21'b101101101000100101000;
		14'b00000111010011:	sigmoid = 21'b101101101010001101110;
		14'b00000111010100:	sigmoid = 21'b101101101011110110011;
		14'b00000111010101:	sigmoid = 21'b101101101101011110111;
		14'b00000111010110:	sigmoid = 21'b101101101111000111011;
		14'b00000111010111:	sigmoid = 21'b101101110000101111110;
		14'b00000111011000:	sigmoid = 21'b101101110010011000000;
		14'b00000111011001:	sigmoid = 21'b101101110100000000010;
		14'b00000111011010:	sigmoid = 21'b101101110101101000011;
		14'b00000111011011:	sigmoid = 21'b101101110111010000011;
		14'b00000111011100:	sigmoid = 21'b101101111000111000010;
		14'b00000111011101:	sigmoid = 21'b101101111010100000001;
		14'b00000111011110:	sigmoid = 21'b101101111100000111111;
		14'b00000111011111:	sigmoid = 21'b101101111101101111101;
		14'b00000111100000:	sigmoid = 21'b101101111111010111001;
		14'b00000111100001:	sigmoid = 21'b101110000000111110101;
		14'b00000111100010:	sigmoid = 21'b101110000010100110000;
		14'b00000111100011:	sigmoid = 21'b101110000100001101011;
		14'b00000111100100:	sigmoid = 21'b101110000101110100101;
		14'b00000111100101:	sigmoid = 21'b101110000111011011110;
		14'b00000111100110:	sigmoid = 21'b101110001001000010110;
		14'b00000111100111:	sigmoid = 21'b101110001010101001110;
		14'b00000111101000:	sigmoid = 21'b101110001100010000101;
		14'b00000111101001:	sigmoid = 21'b101110001101110111011;
		14'b00000111101010:	sigmoid = 21'b101110001111011110000;
		14'b00000111101011:	sigmoid = 21'b101110010001000100101;
		14'b00000111101100:	sigmoid = 21'b101110010010101011001;
		14'b00000111101101:	sigmoid = 21'b101110010100010001101;
		14'b00000111101110:	sigmoid = 21'b101110010101110111111;
		14'b00000111101111:	sigmoid = 21'b101110010111011110001;
		14'b00000111110000:	sigmoid = 21'b101110011001000100011;
		14'b00000111110001:	sigmoid = 21'b101110011010101010011;
		14'b00000111110010:	sigmoid = 21'b101110011100010000011;
		14'b00000111110011:	sigmoid = 21'b101110011101110110010;
		14'b00000111110100:	sigmoid = 21'b101110011111011100000;
		14'b00000111110101:	sigmoid = 21'b101110100001000001110;
		14'b00000111110110:	sigmoid = 21'b101110100010100111011;
		14'b00000111110111:	sigmoid = 21'b101110100100001100111;
		14'b00000111111000:	sigmoid = 21'b101110100101110010011;
		14'b00000111111001:	sigmoid = 21'b101110100111010111101;
		14'b00000111111010:	sigmoid = 21'b101110101000111100111;
		14'b00000111111011:	sigmoid = 21'b101110101010100010001;
		14'b00000111111100:	sigmoid = 21'b101110101100000111001;
		14'b00000111111101:	sigmoid = 21'b101110101101101100001;
		14'b00000111111110:	sigmoid = 21'b101110101111010001000;
		14'b00000111111111:	sigmoid = 21'b101110110000110101111;
		14'b00001000000000:	sigmoid = 21'b101110110010011010100;
		14'b00001000000001:	sigmoid = 21'b101110110011111111001;
		14'b00001000000010:	sigmoid = 21'b101110110101100011110;
		14'b00001000000011:	sigmoid = 21'b101110110111001000001;
		14'b00001000000100:	sigmoid = 21'b101110111000101100100;
		14'b00001000000101:	sigmoid = 21'b101110111010010000110;
		14'b00001000000110:	sigmoid = 21'b101110111011110100111;
		14'b00001000000111:	sigmoid = 21'b101110111101011001000;
		14'b00001000001000:	sigmoid = 21'b101110111110111101000;
		14'b00001000001001:	sigmoid = 21'b101111000000100000111;
		14'b00001000001010:	sigmoid = 21'b101111000010000100101;
		14'b00001000001011:	sigmoid = 21'b101111000011101000011;
		14'b00001000001100:	sigmoid = 21'b101111000101001100000;
		14'b00001000001101:	sigmoid = 21'b101111000110101111100;
		14'b00001000001110:	sigmoid = 21'b101111001000010010111;
		14'b00001000001111:	sigmoid = 21'b101111001001110110010;
		14'b00001000010000:	sigmoid = 21'b101111001011011001100;
		14'b00001000010001:	sigmoid = 21'b101111001100111100101;
		14'b00001000010010:	sigmoid = 21'b101111001110011111110;
		14'b00001000010011:	sigmoid = 21'b101111010000000010110;
		14'b00001000010100:	sigmoid = 21'b101111010001100101101;
		14'b00001000010101:	sigmoid = 21'b101111010011001000011;
		14'b00001000010110:	sigmoid = 21'b101111010100101011001;
		14'b00001000010111:	sigmoid = 21'b101111010110001101110;
		14'b00001000011000:	sigmoid = 21'b101111010111110000010;
		14'b00001000011001:	sigmoid = 21'b101111011001010010101;
		14'b00001000011010:	sigmoid = 21'b101111011010110101000;
		14'b00001000011011:	sigmoid = 21'b101111011100010111001;
		14'b00001000011100:	sigmoid = 21'b101111011101111001011;
		14'b00001000011101:	sigmoid = 21'b101111011111011011011;
		14'b00001000011110:	sigmoid = 21'b101111100000111101011;
		14'b00001000011111:	sigmoid = 21'b101111100010011111010;
		14'b00001000100000:	sigmoid = 21'b101111100100000001000;
		14'b00001000100001:	sigmoid = 21'b101111100101100010101;
		14'b00001000100010:	sigmoid = 21'b101111100111000100010;
		14'b00001000100011:	sigmoid = 21'b101111101000100101110;
		14'b00001000100100:	sigmoid = 21'b101111101010000111001;
		14'b00001000100101:	sigmoid = 21'b101111101011101000011;
		14'b00001000100110:	sigmoid = 21'b101111101101001001101;
		14'b00001000100111:	sigmoid = 21'b101111101110101010110;
		14'b00001000101000:	sigmoid = 21'b101111110000001011110;
		14'b00001000101001:	sigmoid = 21'b101111110001101100110;
		14'b00001000101010:	sigmoid = 21'b101111110011001101101;
		14'b00001000101011:	sigmoid = 21'b101111110100101110011;
		14'b00001000101100:	sigmoid = 21'b101111110110001111000;
		14'b00001000101101:	sigmoid = 21'b101111110111101111100;
		14'b00001000101110:	sigmoid = 21'b101111111001010000000;
		14'b00001000101111:	sigmoid = 21'b101111111010110000011;
		14'b00001000110000:	sigmoid = 21'b101111111100010000101;
		14'b00001000110001:	sigmoid = 21'b101111111101110000111;
		14'b00001000110010:	sigmoid = 21'b101111111111010000111;
		14'b00001000110011:	sigmoid = 21'b110000000000110000111;
		14'b00001000110100:	sigmoid = 21'b110000000010010000111;
		14'b00001000110101:	sigmoid = 21'b110000000011110000101;
		14'b00001000110110:	sigmoid = 21'b110000000101010000011;
		14'b00001000110111:	sigmoid = 21'b110000000110110000000;
		14'b00001000111000:	sigmoid = 21'b110000001000001111100;
		14'b00001000111001:	sigmoid = 21'b110000001001101111000;
		14'b00001000111010:	sigmoid = 21'b110000001011001110010;
		14'b00001000111011:	sigmoid = 21'b110000001100101101100;
		14'b00001000111100:	sigmoid = 21'b110000001110001100110;
		14'b00001000111101:	sigmoid = 21'b110000001111101011110;
		14'b00001000111110:	sigmoid = 21'b110000010001001010110;
		14'b00001000111111:	sigmoid = 21'b110000010010101001101;
		14'b00001001000000:	sigmoid = 21'b110000010100001000011;
		14'b00001001000001:	sigmoid = 21'b110000010101100111000;
		14'b00001001000010:	sigmoid = 21'b110000010111000101101;
		14'b00001001000011:	sigmoid = 21'b110000011000100100001;
		14'b00001001000100:	sigmoid = 21'b110000011010000010100;
		14'b00001001000101:	sigmoid = 21'b110000011011100000111;
		14'b00001001000110:	sigmoid = 21'b110000011100111111000;
		14'b00001001000111:	sigmoid = 21'b110000011110011101001;
		14'b00001001001000:	sigmoid = 21'b110000011111111011001;
		14'b00001001001001:	sigmoid = 21'b110000100001011001001;
		14'b00001001001010:	sigmoid = 21'b110000100010110111000;
		14'b00001001001011:	sigmoid = 21'b110000100100010100101;
		14'b00001001001100:	sigmoid = 21'b110000100101110010011;
		14'b00001001001101:	sigmoid = 21'b110000100111001111111;
		14'b00001001001110:	sigmoid = 21'b110000101000101101011;
		14'b00001001001111:	sigmoid = 21'b110000101010001010101;
		14'b00001001010000:	sigmoid = 21'b110000101011101000000;
		14'b00001001010001:	sigmoid = 21'b110000101101000101001;
		14'b00001001010010:	sigmoid = 21'b110000101110100010001;
		14'b00001001010011:	sigmoid = 21'b110000101111111111001;
		14'b00001001010100:	sigmoid = 21'b110000110001011100000;
		14'b00001001010101:	sigmoid = 21'b110000110010111000111;
		14'b00001001010110:	sigmoid = 21'b110000110100010101100;
		14'b00001001010111:	sigmoid = 21'b110000110101110010001;
		14'b00001001011000:	sigmoid = 21'b110000110111001110101;
		14'b00001001011001:	sigmoid = 21'b110000111000101011000;
		14'b00001001011010:	sigmoid = 21'b110000111010000111011;
		14'b00001001011011:	sigmoid = 21'b110000111011100011100;
		14'b00001001011100:	sigmoid = 21'b110000111100111111101;
		14'b00001001011101:	sigmoid = 21'b110000111110011011110;
		14'b00001001011110:	sigmoid = 21'b110000111111110111101;
		14'b00001001011111:	sigmoid = 21'b110001000001010011100;
		14'b00001001100000:	sigmoid = 21'b110001000010101111010;
		14'b00001001100001:	sigmoid = 21'b110001000100001010111;
		14'b00001001100010:	sigmoid = 21'b110001000101100110011;
		14'b00001001100011:	sigmoid = 21'b110001000111000001111;
		14'b00001001100100:	sigmoid = 21'b110001001000011101010;
		14'b00001001100101:	sigmoid = 21'b110001001001111000100;
		14'b00001001100110:	sigmoid = 21'b110001001011010011101;
		14'b00001001100111:	sigmoid = 21'b110001001100101110110;
		14'b00001001101000:	sigmoid = 21'b110001001110001001110;
		14'b00001001101001:	sigmoid = 21'b110001001111100100101;
		14'b00001001101010:	sigmoid = 21'b110001010000111111011;
		14'b00001001101011:	sigmoid = 21'b110001010010011010001;
		14'b00001001101100:	sigmoid = 21'b110001010011110100101;
		14'b00001001101101:	sigmoid = 21'b110001010101001111001;
		14'b00001001101110:	sigmoid = 21'b110001010110101001100;
		14'b00001001101111:	sigmoid = 21'b110001011000000011111;
		14'b00001001110000:	sigmoid = 21'b110001011001011110001;
		14'b00001001110001:	sigmoid = 21'b110001011010111000010;
		14'b00001001110010:	sigmoid = 21'b110001011100010010010;
		14'b00001001110011:	sigmoid = 21'b110001011101101100001;
		14'b00001001110100:	sigmoid = 21'b110001011111000110000;
		14'b00001001110101:	sigmoid = 21'b110001100000011111110;
		14'b00001001110110:	sigmoid = 21'b110001100001111001011;
		14'b00001001110111:	sigmoid = 21'b110001100011010010111;
		14'b00001001111000:	sigmoid = 21'b110001100100101100011;
		14'b00001001111001:	sigmoid = 21'b110001100110000101101;
		14'b00001001111010:	sigmoid = 21'b110001100111011110111;
		14'b00001001111011:	sigmoid = 21'b110001101000111000001;
		14'b00001001111100:	sigmoid = 21'b110001101010010001001;
		14'b00001001111101:	sigmoid = 21'b110001101011101010001;
		14'b00001001111110:	sigmoid = 21'b110001101101000011000;
		14'b00001001111111:	sigmoid = 21'b110001101110011011110;
		14'b00001010000000:	sigmoid = 21'b110001101111110100011;
		14'b00001010000001:	sigmoid = 21'b110001110001001101000;
		14'b00001010000010:	sigmoid = 21'b110001110010100101100;
		14'b00001010000011:	sigmoid = 21'b110001110011111101111;
		14'b00001010000100:	sigmoid = 21'b110001110101010110001;
		14'b00001010000101:	sigmoid = 21'b110001110110101110011;
		14'b00001010000110:	sigmoid = 21'b110001111000000110100;
		14'b00001010000111:	sigmoid = 21'b110001111001011110100;
		14'b00001010001000:	sigmoid = 21'b110001111010110110011;
		14'b00001010001001:	sigmoid = 21'b110001111100001110010;
		14'b00001010001010:	sigmoid = 21'b110001111101100101111;
		14'b00001010001011:	sigmoid = 21'b110001111110111101100;
		14'b00001010001100:	sigmoid = 21'b110010000000010101001;
		14'b00001010001101:	sigmoid = 21'b110010000001101100100;
		14'b00001010001110:	sigmoid = 21'b110010000011000011111;
		14'b00001010001111:	sigmoid = 21'b110010000100011011001;
		14'b00001010010000:	sigmoid = 21'b110010000101110010010;
		14'b00001010010001:	sigmoid = 21'b110010000111001001010;
		14'b00001010010010:	sigmoid = 21'b110010001000100000010;
		14'b00001010010011:	sigmoid = 21'b110010001001110111000;
		14'b00001010010100:	sigmoid = 21'b110010001011001101110;
		14'b00001010010101:	sigmoid = 21'b110010001100100100100;
		14'b00001010010110:	sigmoid = 21'b110010001101111011000;
		14'b00001010010111:	sigmoid = 21'b110010001111010001100;
		14'b00001010011000:	sigmoid = 21'b110010010000100111111;
		14'b00001010011001:	sigmoid = 21'b110010010001111110001;
		14'b00001010011010:	sigmoid = 21'b110010010011010100011;
		14'b00001010011011:	sigmoid = 21'b110010010100101010011;
		14'b00001010011100:	sigmoid = 21'b110010010110000000011;
		14'b00001010011101:	sigmoid = 21'b110010010111010110010;
		14'b00001010011110:	sigmoid = 21'b110010011000101100001;
		14'b00001010011111:	sigmoid = 21'b110010011010000001110;
		14'b00001010100000:	sigmoid = 21'b110010011011010111011;
		14'b00001010100001:	sigmoid = 21'b110010011100101100111;
		14'b00001010100010:	sigmoid = 21'b110010011110000010010;
		14'b00001010100011:	sigmoid = 21'b110010011111010111101;
		14'b00001010100100:	sigmoid = 21'b110010100000101100111;
		14'b00001010100101:	sigmoid = 21'b110010100010000001111;
		14'b00001010100110:	sigmoid = 21'b110010100011010111000;
		14'b00001010100111:	sigmoid = 21'b110010100100101011111;
		14'b00001010101000:	sigmoid = 21'b110010100110000000110;
		14'b00001010101001:	sigmoid = 21'b110010100111010101100;
		14'b00001010101010:	sigmoid = 21'b110010101000101010001;
		14'b00001010101011:	sigmoid = 21'b110010101001111110101;
		14'b00001010101100:	sigmoid = 21'b110010101011010011001;
		14'b00001010101101:	sigmoid = 21'b110010101100100111011;
		14'b00001010101110:	sigmoid = 21'b110010101101111011101;
		14'b00001010101111:	sigmoid = 21'b110010101111001111111;
		14'b00001010110000:	sigmoid = 21'b110010110000100011111;
		14'b00001010110001:	sigmoid = 21'b110010110001110111111;
		14'b00001010110010:	sigmoid = 21'b110010110011001011110;
		14'b00001010110011:	sigmoid = 21'b110010110100011111100;
		14'b00001010110100:	sigmoid = 21'b110010110101110011010;
		14'b00001010110101:	sigmoid = 21'b110010110111000110110;
		14'b00001010110110:	sigmoid = 21'b110010111000011010010;
		14'b00001010110111:	sigmoid = 21'b110010111001101101101;
		14'b00001010111000:	sigmoid = 21'b110010111011000000111;
		14'b00001010111001:	sigmoid = 21'b110010111100010100001;
		14'b00001010111010:	sigmoid = 21'b110010111101100111010;
		14'b00001010111011:	sigmoid = 21'b110010111110111010010;
		14'b00001010111100:	sigmoid = 21'b110011000000001101001;
		14'b00001010111101:	sigmoid = 21'b110011000001100000000;
		14'b00001010111110:	sigmoid = 21'b110011000010110010101;
		14'b00001010111111:	sigmoid = 21'b110011000100000101010;
		14'b00001011000000:	sigmoid = 21'b110011000101010111110;
		14'b00001011000001:	sigmoid = 21'b110011000110101010010;
		14'b00001011000010:	sigmoid = 21'b110011000111111100101;
		14'b00001011000011:	sigmoid = 21'b110011001001001110110;
		14'b00001011000100:	sigmoid = 21'b110011001010100001000;
		14'b00001011000101:	sigmoid = 21'b110011001011110011000;
		14'b00001011000110:	sigmoid = 21'b110011001101000100111;
		14'b00001011000111:	sigmoid = 21'b110011001110010110110;
		14'b00001011001000:	sigmoid = 21'b110011001111101000100;
		14'b00001011001001:	sigmoid = 21'b110011010000111010010;
		14'b00001011001010:	sigmoid = 21'b110011010010001011110;
		14'b00001011001011:	sigmoid = 21'b110011010011011101010;
		14'b00001011001100:	sigmoid = 21'b110011010100101110101;
		14'b00001011001101:	sigmoid = 21'b110011010101111111111;
		14'b00001011001110:	sigmoid = 21'b110011010111010001000;
		14'b00001011001111:	sigmoid = 21'b110011011000100010001;
		14'b00001011010000:	sigmoid = 21'b110011011001110011001;
		14'b00001011010001:	sigmoid = 21'b110011011011000100000;
		14'b00001011010010:	sigmoid = 21'b110011011100010100111;
		14'b00001011010011:	sigmoid = 21'b110011011101100101100;
		14'b00001011010100:	sigmoid = 21'b110011011110110110001;
		14'b00001011010101:	sigmoid = 21'b110011100000000110101;
		14'b00001011010110:	sigmoid = 21'b110011100001010111000;
		14'b00001011010111:	sigmoid = 21'b110011100010100111011;
		14'b00001011011000:	sigmoid = 21'b110011100011110111101;
		14'b00001011011001:	sigmoid = 21'b110011100101000111110;
		14'b00001011011010:	sigmoid = 21'b110011100110010111110;
		14'b00001011011011:	sigmoid = 21'b110011100111100111101;
		14'b00001011011100:	sigmoid = 21'b110011101000110111100;
		14'b00001011011101:	sigmoid = 21'b110011101010000111010;
		14'b00001011011110:	sigmoid = 21'b110011101011010110111;
		14'b00001011011111:	sigmoid = 21'b110011101100100110100;
		14'b00001011100000:	sigmoid = 21'b110011101101110101111;
		14'b00001011100001:	sigmoid = 21'b110011101111000101010;
		14'b00001011100010:	sigmoid = 21'b110011110000010100100;
		14'b00001011100011:	sigmoid = 21'b110011110001100011110;
		14'b00001011100100:	sigmoid = 21'b110011110010110010110;
		14'b00001011100101:	sigmoid = 21'b110011110100000001110;
		14'b00001011100110:	sigmoid = 21'b110011110101010000101;
		14'b00001011100111:	sigmoid = 21'b110011110110011111011;
		14'b00001011101000:	sigmoid = 21'b110011110111101110001;
		14'b00001011101001:	sigmoid = 21'b110011111000111100110;
		14'b00001011101010:	sigmoid = 21'b110011111010001011010;
		14'b00001011101011:	sigmoid = 21'b110011111011011001101;
		14'b00001011101100:	sigmoid = 21'b110011111100100111111;
		14'b00001011101101:	sigmoid = 21'b110011111101110110001;
		14'b00001011101110:	sigmoid = 21'b110011111111000100010;
		14'b00001011101111:	sigmoid = 21'b110100000000010010010;
		14'b00001011110000:	sigmoid = 21'b110100000001100000010;
		14'b00001011110001:	sigmoid = 21'b110100000010101110000;
		14'b00001011110010:	sigmoid = 21'b110100000011111011110;
		14'b00001011110011:	sigmoid = 21'b110100000101001001100;
		14'b00001011110100:	sigmoid = 21'b110100000110010111000;
		14'b00001011110101:	sigmoid = 21'b110100000111100100100;
		14'b00001011110110:	sigmoid = 21'b110100001000110001110;
		14'b00001011110111:	sigmoid = 21'b110100001001111111001;
		14'b00001011111000:	sigmoid = 21'b110100001011001100010;
		14'b00001011111001:	sigmoid = 21'b110100001100011001011;
		14'b00001011111010:	sigmoid = 21'b110100001101100110010;
		14'b00001011111011:	sigmoid = 21'b110100001110110011001;
		14'b00001011111100:	sigmoid = 21'b110100010000000000000;
		14'b00001011111101:	sigmoid = 21'b110100010001001100101;
		14'b00001011111110:	sigmoid = 21'b110100010010011001010;
		14'b00001011111111:	sigmoid = 21'b110100010011100101110;
		14'b00001100000000:	sigmoid = 21'b110100010100110010001;
		14'b00001100000001:	sigmoid = 21'b110100010101111110100;
		14'b00001100000010:	sigmoid = 21'b110100010111001010110;
		14'b00001100000011:	sigmoid = 21'b110100011000010110111;
		14'b00001100000100:	sigmoid = 21'b110100011001100010111;
		14'b00001100000101:	sigmoid = 21'b110100011010101110110;
		14'b00001100000110:	sigmoid = 21'b110100011011111010101;
		14'b00001100000111:	sigmoid = 21'b110100011101000110011;
		14'b00001100001000:	sigmoid = 21'b110100011110010010000;
		14'b00001100001001:	sigmoid = 21'b110100011111011101101;
		14'b00001100001010:	sigmoid = 21'b110100100000101001001;
		14'b00001100001011:	sigmoid = 21'b110100100001110100100;
		14'b00001100001100:	sigmoid = 21'b110100100010111111110;
		14'b00001100001101:	sigmoid = 21'b110100100100001010111;
		14'b00001100001110:	sigmoid = 21'b110100100101010110000;
		14'b00001100001111:	sigmoid = 21'b110100100110100001000;
		14'b00001100010000:	sigmoid = 21'b110100100111101011111;
		14'b00001100010001:	sigmoid = 21'b110100101000110110110;
		14'b00001100010010:	sigmoid = 21'b110100101010000001011;
		14'b00001100010011:	sigmoid = 21'b110100101011001100000;
		14'b00001100010100:	sigmoid = 21'b110100101100010110100;
		14'b00001100010101:	sigmoid = 21'b110100101101100001000;
		14'b00001100010110:	sigmoid = 21'b110100101110101011010;
		14'b00001100010111:	sigmoid = 21'b110100101111110101100;
		14'b00001100011000:	sigmoid = 21'b110100110000111111101;
		14'b00001100011001:	sigmoid = 21'b110100110010001001110;
		14'b00001100011010:	sigmoid = 21'b110100110011010011110;
		14'b00001100011011:	sigmoid = 21'b110100110100011101100;
		14'b00001100011100:	sigmoid = 21'b110100110101100111011;
		14'b00001100011101:	sigmoid = 21'b110100110110110001000;
		14'b00001100011110:	sigmoid = 21'b110100110111111010101;
		14'b00001100011111:	sigmoid = 21'b110100111001000100001;
		14'b00001100100000:	sigmoid = 21'b110100111010001101100;
		14'b00001100100001:	sigmoid = 21'b110100111011010110110;
		14'b00001100100010:	sigmoid = 21'b110100111100100000000;
		14'b00001100100011:	sigmoid = 21'b110100111101101001001;
		14'b00001100100100:	sigmoid = 21'b110100111110110010001;
		14'b00001100100101:	sigmoid = 21'b110100111111111011000;
		14'b00001100100110:	sigmoid = 21'b110101000001000011111;
		14'b00001100100111:	sigmoid = 21'b110101000010001100101;
		14'b00001100101000:	sigmoid = 21'b110101000011010101010;
		14'b00001100101001:	sigmoid = 21'b110101000100011101111;
		14'b00001100101010:	sigmoid = 21'b110101000101100110010;
		14'b00001100101011:	sigmoid = 21'b110101000110101110101;
		14'b00001100101100:	sigmoid = 21'b110101000111110110111;
		14'b00001100101101:	sigmoid = 21'b110101001000111111001;
		14'b00001100101110:	sigmoid = 21'b110101001010000111010;
		14'b00001100101111:	sigmoid = 21'b110101001011001111010;
		14'b00001100110000:	sigmoid = 21'b110101001100010111001;
		14'b00001100110001:	sigmoid = 21'b110101001101011110111;
		14'b00001100110010:	sigmoid = 21'b110101001110100110101;
		14'b00001100110011:	sigmoid = 21'b110101001111101110010;
		14'b00001100110100:	sigmoid = 21'b110101010000110101110;
		14'b00001100110101:	sigmoid = 21'b110101010001111101010;
		14'b00001100110110:	sigmoid = 21'b110101010011000100101;
		14'b00001100110111:	sigmoid = 21'b110101010100001011111;
		14'b00001100111000:	sigmoid = 21'b110101010101010011000;
		14'b00001100111001:	sigmoid = 21'b110101010110011010000;
		14'b00001100111010:	sigmoid = 21'b110101010111100001000;
		14'b00001100111011:	sigmoid = 21'b110101011000100111111;
		14'b00001100111100:	sigmoid = 21'b110101011001101110110;
		14'b00001100111101:	sigmoid = 21'b110101011010110101011;
		14'b00001100111110:	sigmoid = 21'b110101011011111100000;
		14'b00001100111111:	sigmoid = 21'b110101011101000010100;
		14'b00001101000000:	sigmoid = 21'b110101011110001000111;
		14'b00001101000001:	sigmoid = 21'b110101011111001111010;
		14'b00001101000010:	sigmoid = 21'b110101100000010101100;
		14'b00001101000011:	sigmoid = 21'b110101100001011011101;
		14'b00001101000100:	sigmoid = 21'b110101100010100001110;
		14'b00001101000101:	sigmoid = 21'b110101100011100111101;
		14'b00001101000110:	sigmoid = 21'b110101100100101101100;
		14'b00001101000111:	sigmoid = 21'b110101100101110011010;
		14'b00001101001000:	sigmoid = 21'b110101100110111001000;
		14'b00001101001001:	sigmoid = 21'b110101100111111110101;
		14'b00001101001010:	sigmoid = 21'b110101101001000100001;
		14'b00001101001011:	sigmoid = 21'b110101101010001001100;
		14'b00001101001100:	sigmoid = 21'b110101101011001110110;
		14'b00001101001101:	sigmoid = 21'b110101101100010100000;
		14'b00001101001110:	sigmoid = 21'b110101101101011001001;
		14'b00001101001111:	sigmoid = 21'b110101101110011110010;
		14'b00001101010000:	sigmoid = 21'b110101101111100011001;
		14'b00001101010001:	sigmoid = 21'b110101110000101000000;
		14'b00001101010010:	sigmoid = 21'b110101110001101100110;
		14'b00001101010011:	sigmoid = 21'b110101110010110001100;
		14'b00001101010100:	sigmoid = 21'b110101110011110110000;
		14'b00001101010101:	sigmoid = 21'b110101110100111010100;
		14'b00001101010110:	sigmoid = 21'b110101110101111111000;
		14'b00001101010111:	sigmoid = 21'b110101110111000011010;
		14'b00001101011000:	sigmoid = 21'b110101111000000111100;
		14'b00001101011001:	sigmoid = 21'b110101111001001011101;
		14'b00001101011010:	sigmoid = 21'b110101111010001111101;
		14'b00001101011011:	sigmoid = 21'b110101111011010011101;
		14'b00001101011100:	sigmoid = 21'b110101111100010111100;
		14'b00001101011101:	sigmoid = 21'b110101111101011011010;
		14'b00001101011110:	sigmoid = 21'b110101111110011110111;
		14'b00001101011111:	sigmoid = 21'b110101111111100010100;
		14'b00001101100000:	sigmoid = 21'b110110000000100110000;
		14'b00001101100001:	sigmoid = 21'b110110000001101001011;
		14'b00001101100010:	sigmoid = 21'b110110000010101100110;
		14'b00001101100011:	sigmoid = 21'b110110000011101111111;
		14'b00001101100100:	sigmoid = 21'b110110000100110011000;
		14'b00001101100101:	sigmoid = 21'b110110000101110110001;
		14'b00001101100110:	sigmoid = 21'b110110000110111001000;
		14'b00001101100111:	sigmoid = 21'b110110000111111011111;
		14'b00001101101000:	sigmoid = 21'b110110001000111110101;
		14'b00001101101001:	sigmoid = 21'b110110001010000001011;
		14'b00001101101010:	sigmoid = 21'b110110001011000100000;
		14'b00001101101011:	sigmoid = 21'b110110001100000110100;
		14'b00001101101100:	sigmoid = 21'b110110001101001000111;
		14'b00001101101101:	sigmoid = 21'b110110001110001011001;
		14'b00001101101110:	sigmoid = 21'b110110001111001101011;
		14'b00001101101111:	sigmoid = 21'b110110010000001111100;
		14'b00001101110000:	sigmoid = 21'b110110010001010001101;
		14'b00001101110001:	sigmoid = 21'b110110010010010011100;
		14'b00001101110010:	sigmoid = 21'b110110010011010101011;
		14'b00001101110011:	sigmoid = 21'b110110010100010111010;
		14'b00001101110100:	sigmoid = 21'b110110010101011000111;
		14'b00001101110101:	sigmoid = 21'b110110010110011010100;
		14'b00001101110110:	sigmoid = 21'b110110010111011100000;
		14'b00001101110111:	sigmoid = 21'b110110011000011101100;
		14'b00001101111000:	sigmoid = 21'b110110011001011110110;
		14'b00001101111001:	sigmoid = 21'b110110011010100000000;
		14'b00001101111010:	sigmoid = 21'b110110011011100001001;
		14'b00001101111011:	sigmoid = 21'b110110011100100010010;
		14'b00001101111100:	sigmoid = 21'b110110011101100011010;
		14'b00001101111101:	sigmoid = 21'b110110011110100100001;
		14'b00001101111110:	sigmoid = 21'b110110011111100100111;
		14'b00001101111111:	sigmoid = 21'b110110100000100101101;
		14'b00001110000000:	sigmoid = 21'b110110100001100110010;
		14'b00001110000001:	sigmoid = 21'b110110100010100110110;
		14'b00001110000010:	sigmoid = 21'b110110100011100111010;
		14'b00001110000011:	sigmoid = 21'b110110100100100111101;
		14'b00001110000100:	sigmoid = 21'b110110100101100111111;
		14'b00001110000101:	sigmoid = 21'b110110100110101000000;
		14'b00001110000110:	sigmoid = 21'b110110100111101000001;
		14'b00001110000111:	sigmoid = 21'b110110101000101000001;
		14'b00001110001000:	sigmoid = 21'b110110101001101000000;
		14'b00001110001001:	sigmoid = 21'b110110101010100111111;
		14'b00001110001010:	sigmoid = 21'b110110101011100111101;
		14'b00001110001011:	sigmoid = 21'b110110101100100111010;
		14'b00001110001100:	sigmoid = 21'b110110101101100110111;
		14'b00001110001101:	sigmoid = 21'b110110101110100110010;
		14'b00001110001110:	sigmoid = 21'b110110101111100101101;
		14'b00001110001111:	sigmoid = 21'b110110110000100101000;
		14'b00001110010000:	sigmoid = 21'b110110110001100100001;
		14'b00001110010001:	sigmoid = 21'b110110110010100011010;
		14'b00001110010010:	sigmoid = 21'b110110110011100010011;
		14'b00001110010011:	sigmoid = 21'b110110110100100001010;
		14'b00001110010100:	sigmoid = 21'b110110110101100000001;
		14'b00001110010101:	sigmoid = 21'b110110110110011110111;
		14'b00001110010110:	sigmoid = 21'b110110110111011101101;
		14'b00001110010111:	sigmoid = 21'b110110111000011100010;
		14'b00001110011000:	sigmoid = 21'b110110111001011010110;
		14'b00001110011001:	sigmoid = 21'b110110111010011001001;
		14'b00001110011010:	sigmoid = 21'b110110111011010111100;
		14'b00001110011011:	sigmoid = 21'b110110111100010101110;
		14'b00001110011100:	sigmoid = 21'b110110111101010011111;
		14'b00001110011101:	sigmoid = 21'b110110111110010001111;
		14'b00001110011110:	sigmoid = 21'b110110111111001111111;
		14'b00001110011111:	sigmoid = 21'b110111000000001101111;
		14'b00001110100000:	sigmoid = 21'b110111000001001011101;
		14'b00001110100001:	sigmoid = 21'b110111000010001001011;
		14'b00001110100010:	sigmoid = 21'b110111000011000111000;
		14'b00001110100011:	sigmoid = 21'b110111000100000100100;
		14'b00001110100100:	sigmoid = 21'b110111000101000010000;
		14'b00001110100101:	sigmoid = 21'b110111000101111111011;
		14'b00001110100110:	sigmoid = 21'b110111000110111100101;
		14'b00001110100111:	sigmoid = 21'b110111000111111001111;
		14'b00001110101000:	sigmoid = 21'b110111001000110111000;
		14'b00001110101001:	sigmoid = 21'b110111001001110100000;
		14'b00001110101010:	sigmoid = 21'b110111001010110001000;
		14'b00001110101011:	sigmoid = 21'b110111001011101101111;
		14'b00001110101100:	sigmoid = 21'b110111001100101010101;
		14'b00001110101101:	sigmoid = 21'b110111001101100111011;
		14'b00001110101110:	sigmoid = 21'b110111001110100011111;
		14'b00001110101111:	sigmoid = 21'b110111001111100000011;
		14'b00001110110000:	sigmoid = 21'b110111010000011100111;
		14'b00001110110001:	sigmoid = 21'b110111010001011001010;
		14'b00001110110010:	sigmoid = 21'b110111010010010101100;
		14'b00001110110011:	sigmoid = 21'b110111010011010001101;
		14'b00001110110100:	sigmoid = 21'b110111010100001101110;
		14'b00001110110101:	sigmoid = 21'b110111010101001001110;
		14'b00001110110110:	sigmoid = 21'b110111010110000101101;
		14'b00001110110111:	sigmoid = 21'b110111010111000001100;
		14'b00001110111000:	sigmoid = 21'b110111010111111101010;
		14'b00001110111001:	sigmoid = 21'b110111011000111000111;
		14'b00001110111010:	sigmoid = 21'b110111011001110100100;
		14'b00001110111011:	sigmoid = 21'b110111011010110000000;
		14'b00001110111100:	sigmoid = 21'b110111011011101011011;
		14'b00001110111101:	sigmoid = 21'b110111011100100110110;
		14'b00001110111110:	sigmoid = 21'b110111011101100010000;
		14'b00001110111111:	sigmoid = 21'b110111011110011101001;
		14'b00001111000000:	sigmoid = 21'b110111011111011000001;
		14'b00001111000001:	sigmoid = 21'b110111100000010011001;
		14'b00001111000010:	sigmoid = 21'b110111100001001110000;
		14'b00001111000011:	sigmoid = 21'b110111100010001000111;
		14'b00001111000100:	sigmoid = 21'b110111100011000011101;
		14'b00001111000101:	sigmoid = 21'b110111100011111110010;
		14'b00001111000110:	sigmoid = 21'b110111100100111000110;
		14'b00001111000111:	sigmoid = 21'b110111100101110011010;
		14'b00001111001000:	sigmoid = 21'b110111100110101101101;
		14'b00001111001001:	sigmoid = 21'b110111100111101000000;
		14'b00001111001010:	sigmoid = 21'b110111101000100010010;
		14'b00001111001011:	sigmoid = 21'b110111101001011100011;
		14'b00001111001100:	sigmoid = 21'b110111101010010110011;
		14'b00001111001101:	sigmoid = 21'b110111101011010000011;
		14'b00001111001110:	sigmoid = 21'b110111101100001010010;
		14'b00001111001111:	sigmoid = 21'b110111101101000100001;
		14'b00001111010000:	sigmoid = 21'b110111101101111101110;
		14'b00001111010001:	sigmoid = 21'b110111101110110111011;
		14'b00001111010010:	sigmoid = 21'b110111101111110001000;
		14'b00001111010011:	sigmoid = 21'b110111110000101010100;
		14'b00001111010100:	sigmoid = 21'b110111110001100011111;
		14'b00001111010101:	sigmoid = 21'b110111110010011101001;
		14'b00001111010110:	sigmoid = 21'b110111110011010110011;
		14'b00001111010111:	sigmoid = 21'b110111110100001111100;
		14'b00001111011000:	sigmoid = 21'b110111110101001000101;
		14'b00001111011001:	sigmoid = 21'b110111110110000001100;
		14'b00001111011010:	sigmoid = 21'b110111110110111010011;
		14'b00001111011011:	sigmoid = 21'b110111110111110011010;
		14'b00001111011100:	sigmoid = 21'b110111111000101100000;
		14'b00001111011101:	sigmoid = 21'b110111111001100100101;
		14'b00001111011110:	sigmoid = 21'b110111111010011101001;
		14'b00001111011111:	sigmoid = 21'b110111111011010101101;
		14'b00001111100000:	sigmoid = 21'b110111111100001110000;
		14'b00001111100001:	sigmoid = 21'b110111111101000110011;
		14'b00001111100010:	sigmoid = 21'b110111111101111110101;
		14'b00001111100011:	sigmoid = 21'b110111111110110110110;
		14'b00001111100100:	sigmoid = 21'b110111111111101110110;
		14'b00001111100101:	sigmoid = 21'b111000000000100110110;
		14'b00001111100110:	sigmoid = 21'b111000000001011110101;
		14'b00001111100111:	sigmoid = 21'b111000000010010110100;
		14'b00001111101000:	sigmoid = 21'b111000000011001110010;
		14'b00001111101001:	sigmoid = 21'b111000000100000101111;
		14'b00001111101010:	sigmoid = 21'b111000000100111101100;
		14'b00001111101011:	sigmoid = 21'b111000000101110101000;
		14'b00001111101100:	sigmoid = 21'b111000000110101100011;
		14'b00001111101101:	sigmoid = 21'b111000000111100011110;
		14'b00001111101110:	sigmoid = 21'b111000001000011011000;
		14'b00001111101111:	sigmoid = 21'b111000001001010010001;
		14'b00001111110000:	sigmoid = 21'b111000001010001001010;
		14'b00001111110001:	sigmoid = 21'b111000001011000000010;
		14'b00001111110010:	sigmoid = 21'b111000001011110111001;
		14'b00001111110011:	sigmoid = 21'b111000001100101110000;
		14'b00001111110100:	sigmoid = 21'b111000001101100100110;
		14'b00001111110101:	sigmoid = 21'b111000001110011011011;
		14'b00001111110110:	sigmoid = 21'b111000001111010010000;
		14'b00001111110111:	sigmoid = 21'b111000010000001000100;
		14'b00001111111000:	sigmoid = 21'b111000010000111111000;
		14'b00001111111001:	sigmoid = 21'b111000010001110101011;
		14'b00001111111010:	sigmoid = 21'b111000010010101011101;
		14'b00001111111011:	sigmoid = 21'b111000010011100001111;
		14'b00001111111100:	sigmoid = 21'b111000010100011000000;
		14'b00001111111101:	sigmoid = 21'b111000010101001110000;
		14'b00001111111110:	sigmoid = 21'b111000010110000011111;
		14'b00001111111111:	sigmoid = 21'b111000010110111001110;
		14'b00010000000000:	sigmoid = 21'b111000010111101111101;
		14'b00010000000001:	sigmoid = 21'b111000011000100101011;
		14'b00010000000010:	sigmoid = 21'b111000011001011011000;
		14'b00010000000011:	sigmoid = 21'b111000011010010000100;
		14'b00010000000100:	sigmoid = 21'b111000011011000110000;
		14'b00010000000101:	sigmoid = 21'b111000011011111011011;
		14'b00010000000110:	sigmoid = 21'b111000011100110000110;
		14'b00010000000111:	sigmoid = 21'b111000011101100110000;
		14'b00010000001000:	sigmoid = 21'b111000011110011011001;
		14'b00010000001001:	sigmoid = 21'b111000011111010000010;
		14'b00010000001010:	sigmoid = 21'b111000100000000101010;
		14'b00010000001011:	sigmoid = 21'b111000100000111010001;
		14'b00010000001100:	sigmoid = 21'b111000100001101111000;
		14'b00010000001101:	sigmoid = 21'b111000100010100011110;
		14'b00010000001110:	sigmoid = 21'b111000100011011000011;
		14'b00010000001111:	sigmoid = 21'b111000100100001101000;
		14'b00010000010000:	sigmoid = 21'b111000100101000001100;
		14'b00010000010001:	sigmoid = 21'b111000100101110110000;
		14'b00010000010010:	sigmoid = 21'b111000100110101010011;
		14'b00010000010011:	sigmoid = 21'b111000100111011110101;
		14'b00010000010100:	sigmoid = 21'b111000101000010010111;
		14'b00010000010101:	sigmoid = 21'b111000101001000111000;
		14'b00010000010110:	sigmoid = 21'b111000101001111011000;
		14'b00010000010111:	sigmoid = 21'b111000101010101111000;
		14'b00010000011000:	sigmoid = 21'b111000101011100010111;
		14'b00010000011001:	sigmoid = 21'b111000101100010110110;
		14'b00010000011010:	sigmoid = 21'b111000101101001010100;
		14'b00010000011011:	sigmoid = 21'b111000101101111110001;
		14'b00010000011100:	sigmoid = 21'b111000101110110001110;
		14'b00010000011101:	sigmoid = 21'b111000101111100101010;
		14'b00010000011110:	sigmoid = 21'b111000110000011000101;
		14'b00010000011111:	sigmoid = 21'b111000110001001100000;
		14'b00010000100000:	sigmoid = 21'b111000110001111111010;
		14'b00010000100001:	sigmoid = 21'b111000110010110010100;
		14'b00010000100010:	sigmoid = 21'b111000110011100101101;
		14'b00010000100011:	sigmoid = 21'b111000110100011000101;
		14'b00010000100100:	sigmoid = 21'b111000110101001011101;
		14'b00010000100101:	sigmoid = 21'b111000110101111110100;
		14'b00010000100110:	sigmoid = 21'b111000110110110001011;
		14'b00010000100111:	sigmoid = 21'b111000110111100100001;
		14'b00010000101000:	sigmoid = 21'b111000111000010110110;
		14'b00010000101001:	sigmoid = 21'b111000111001001001010;
		14'b00010000101010:	sigmoid = 21'b111000111001111011110;
		14'b00010000101011:	sigmoid = 21'b111000111010101110010;
		14'b00010000101100:	sigmoid = 21'b111000111011100000101;
		14'b00010000101101:	sigmoid = 21'b111000111100010010111;
		14'b00010000101110:	sigmoid = 21'b111000111101000101000;
		14'b00010000101111:	sigmoid = 21'b111000111101110111001;
		14'b00010000110000:	sigmoid = 21'b111000111110101001010;
		14'b00010000110001:	sigmoid = 21'b111000111111011011010;
		14'b00010000110010:	sigmoid = 21'b111001000000001101001;
		14'b00010000110011:	sigmoid = 21'b111001000000111110111;
		14'b00010000110100:	sigmoid = 21'b111001000001110000101;
		14'b00010000110101:	sigmoid = 21'b111001000010100010010;
		14'b00010000110110:	sigmoid = 21'b111001000011010011111;
		14'b00010000110111:	sigmoid = 21'b111001000100000101011;
		14'b00010000111000:	sigmoid = 21'b111001000100110110111;
		14'b00010000111001:	sigmoid = 21'b111001000101101000010;
		14'b00010000111010:	sigmoid = 21'b111001000110011001100;
		14'b00010000111011:	sigmoid = 21'b111001000111001010110;
		14'b00010000111100:	sigmoid = 21'b111001000111111011111;
		14'b00010000111101:	sigmoid = 21'b111001001000101100111;
		14'b00010000111110:	sigmoid = 21'b111001001001011101111;
		14'b00010000111111:	sigmoid = 21'b111001001010001110110;
		14'b00010001000000:	sigmoid = 21'b111001001010111111101;
		14'b00010001000001:	sigmoid = 21'b111001001011110000011;
		14'b00010001000010:	sigmoid = 21'b111001001100100001001;
		14'b00010001000011:	sigmoid = 21'b111001001101010001110;
		14'b00010001000100:	sigmoid = 21'b111001001110000010010;
		14'b00010001000101:	sigmoid = 21'b111001001110110010110;
		14'b00010001000110:	sigmoid = 21'b111001001111100011001;
		14'b00010001000111:	sigmoid = 21'b111001010000010011011;
		14'b00010001001000:	sigmoid = 21'b111001010001000011101;
		14'b00010001001001:	sigmoid = 21'b111001010001110011110;
		14'b00010001001010:	sigmoid = 21'b111001010010100011111;
		14'b00010001001011:	sigmoid = 21'b111001010011010011111;
		14'b00010001001100:	sigmoid = 21'b111001010100000011111;
		14'b00010001001101:	sigmoid = 21'b111001010100110011110;
		14'b00010001001110:	sigmoid = 21'b111001010101100011100;
		14'b00010001001111:	sigmoid = 21'b111001010110010011010;
		14'b00010001010000:	sigmoid = 21'b111001010111000010111;
		14'b00010001010001:	sigmoid = 21'b111001010111110010011;
		14'b00010001010010:	sigmoid = 21'b111001011000100001111;
		14'b00010001010011:	sigmoid = 21'b111001011001010001011;
		14'b00010001010100:	sigmoid = 21'b111001011010000000110;
		14'b00010001010101:	sigmoid = 21'b111001011010110000000;
		14'b00010001010110:	sigmoid = 21'b111001011011011111001;
		14'b00010001010111:	sigmoid = 21'b111001011100001110011;
		14'b00010001011000:	sigmoid = 21'b111001011100111101011;
		14'b00010001011001:	sigmoid = 21'b111001011101101100011;
		14'b00010001011010:	sigmoid = 21'b111001011110011011010;
		14'b00010001011011:	sigmoid = 21'b111001011111001010001;
		14'b00010001011100:	sigmoid = 21'b111001011111111000111;
		14'b00010001011101:	sigmoid = 21'b111001100000100111101;
		14'b00010001011110:	sigmoid = 21'b111001100001010110010;
		14'b00010001011111:	sigmoid = 21'b111001100010000100110;
		14'b00010001100000:	sigmoid = 21'b111001100010110011010;
		14'b00010001100001:	sigmoid = 21'b111001100011100001101;
		14'b00010001100010:	sigmoid = 21'b111001100100010000000;
		14'b00010001100011:	sigmoid = 21'b111001100100111110010;
		14'b00010001100100:	sigmoid = 21'b111001100101101100011;
		14'b00010001100101:	sigmoid = 21'b111001100110011010100;
		14'b00010001100110:	sigmoid = 21'b111001100111001000100;
		14'b00010001100111:	sigmoid = 21'b111001100111110110100;
		14'b00010001101000:	sigmoid = 21'b111001101000100100011;
		14'b00010001101001:	sigmoid = 21'b111001101001010010010;
		14'b00010001101010:	sigmoid = 21'b111001101010000000000;
		14'b00010001101011:	sigmoid = 21'b111001101010101101101;
		14'b00010001101100:	sigmoid = 21'b111001101011011011010;
		14'b00010001101101:	sigmoid = 21'b111001101100001000111;
		14'b00010001101110:	sigmoid = 21'b111001101100110110010;
		14'b00010001101111:	sigmoid = 21'b111001101101100011110;
		14'b00010001110000:	sigmoid = 21'b111001101110010001000;
		14'b00010001110001:	sigmoid = 21'b111001101110111110010;
		14'b00010001110010:	sigmoid = 21'b111001101111101011100;
		14'b00010001110011:	sigmoid = 21'b111001110000011000101;
		14'b00010001110100:	sigmoid = 21'b111001110001000101101;
		14'b00010001110101:	sigmoid = 21'b111001110001110010101;
		14'b00010001110110:	sigmoid = 21'b111001110010011111100;
		14'b00010001110111:	sigmoid = 21'b111001110011001100011;
		14'b00010001111000:	sigmoid = 21'b111001110011111001001;
		14'b00010001111001:	sigmoid = 21'b111001110100100101110;
		14'b00010001111010:	sigmoid = 21'b111001110101010010011;
		14'b00010001111011:	sigmoid = 21'b111001110101111111000;
		14'b00010001111100:	sigmoid = 21'b111001110110101011011;
		14'b00010001111101:	sigmoid = 21'b111001110111010111111;
		14'b00010001111110:	sigmoid = 21'b111001111000000100001;
		14'b00010001111111:	sigmoid = 21'b111001111000110000100;
		14'b00010010000000:	sigmoid = 21'b111001111001011100101;
		14'b00010010000001:	sigmoid = 21'b111001111010001000110;
		14'b00010010000010:	sigmoid = 21'b111001111010110100111;
		14'b00010010000011:	sigmoid = 21'b111001111011100000111;
		14'b00010010000100:	sigmoid = 21'b111001111100001100110;
		14'b00010010000101:	sigmoid = 21'b111001111100111000101;
		14'b00010010000110:	sigmoid = 21'b111001111101100100011;
		14'b00010010000111:	sigmoid = 21'b111001111110010000001;
		14'b00010010001000:	sigmoid = 21'b111001111110111011110;
		14'b00010010001001:	sigmoid = 21'b111001111111100111010;
		14'b00010010001010:	sigmoid = 21'b111010000000010010110;
		14'b00010010001011:	sigmoid = 21'b111010000000111110010;
		14'b00010010001100:	sigmoid = 21'b111010000001101001101;
		14'b00010010001101:	sigmoid = 21'b111010000010010100111;
		14'b00010010001110:	sigmoid = 21'b111010000011000000001;
		14'b00010010001111:	sigmoid = 21'b111010000011101011010;
		14'b00010010010000:	sigmoid = 21'b111010000100010110011;
		14'b00010010010001:	sigmoid = 21'b111010000101000001011;
		14'b00010010010010:	sigmoid = 21'b111010000101101100011;
		14'b00010010010011:	sigmoid = 21'b111010000110010111010;
		14'b00010010010100:	sigmoid = 21'b111010000111000010001;
		14'b00010010010101:	sigmoid = 21'b111010000111101100111;
		14'b00010010010110:	sigmoid = 21'b111010001000010111100;
		14'b00010010010111:	sigmoid = 21'b111010001001000010001;
		14'b00010010011000:	sigmoid = 21'b111010001001101100101;
		14'b00010010011001:	sigmoid = 21'b111010001010010111001;
		14'b00010010011010:	sigmoid = 21'b111010001011000001100;
		14'b00010010011011:	sigmoid = 21'b111010001011101011111;
		14'b00010010011100:	sigmoid = 21'b111010001100010110001;
		14'b00010010011101:	sigmoid = 21'b111010001101000000011;
		14'b00010010011110:	sigmoid = 21'b111010001101101010100;
		14'b00010010011111:	sigmoid = 21'b111010001110010100101;
		14'b00010010100000:	sigmoid = 21'b111010001110111110101;
		14'b00010010100001:	sigmoid = 21'b111010001111101000100;
		14'b00010010100010:	sigmoid = 21'b111010010000010010011;
		14'b00010010100011:	sigmoid = 21'b111010010000111100010;
		14'b00010010100100:	sigmoid = 21'b111010010001100110000;
		14'b00010010100101:	sigmoid = 21'b111010010010001111101;
		14'b00010010100110:	sigmoid = 21'b111010010010111001010;
		14'b00010010100111:	sigmoid = 21'b111010010011100010110;
		14'b00010010101000:	sigmoid = 21'b111010010100001100010;
		14'b00010010101001:	sigmoid = 21'b111010010100110101101;
		14'b00010010101010:	sigmoid = 21'b111010010101011111000;
		14'b00010010101011:	sigmoid = 21'b111010010110001000010;
		14'b00010010101100:	sigmoid = 21'b111010010110110001100;
		14'b00010010101101:	sigmoid = 21'b111010010111011010101;
		14'b00010010101110:	sigmoid = 21'b111010011000000011101;
		14'b00010010101111:	sigmoid = 21'b111010011000101100101;
		14'b00010010110000:	sigmoid = 21'b111010011001010101101;
		14'b00010010110001:	sigmoid = 21'b111010011001111110100;
		14'b00010010110010:	sigmoid = 21'b111010011010100111010;
		14'b00010010110011:	sigmoid = 21'b111010011011010000000;
		14'b00010010110100:	sigmoid = 21'b111010011011111000110;
		14'b00010010110101:	sigmoid = 21'b111010011100100001011;
		14'b00010010110110:	sigmoid = 21'b111010011101001001111;
		14'b00010010110111:	sigmoid = 21'b111010011101110010011;
		14'b00010010111000:	sigmoid = 21'b111010011110011010110;
		14'b00010010111001:	sigmoid = 21'b111010011111000011001;
		14'b00010010111010:	sigmoid = 21'b111010011111101011011;
		14'b00010010111011:	sigmoid = 21'b111010100000010011101;
		14'b00010010111100:	sigmoid = 21'b111010100000111011110;
		14'b00010010111101:	sigmoid = 21'b111010100001100011111;
		14'b00010010111110:	sigmoid = 21'b111010100010001011111;
		14'b00010010111111:	sigmoid = 21'b111010100010110011111;
		14'b00010011000000:	sigmoid = 21'b111010100011011011110;
		14'b00010011000001:	sigmoid = 21'b111010100100000011101;
		14'b00010011000010:	sigmoid = 21'b111010100100101011011;
		14'b00010011000011:	sigmoid = 21'b111010100101010011000;
		14'b00010011000100:	sigmoid = 21'b111010100101111010101;
		14'b00010011000101:	sigmoid = 21'b111010100110100010010;
		14'b00010011000110:	sigmoid = 21'b111010100111001001110;
		14'b00010011000111:	sigmoid = 21'b111010100111110001010;
		14'b00010011001000:	sigmoid = 21'b111010101000011000101;
		14'b00010011001001:	sigmoid = 21'b111010101000111111111;
		14'b00010011001010:	sigmoid = 21'b111010101001100111001;
		14'b00010011001011:	sigmoid = 21'b111010101010001110011;
		14'b00010011001100:	sigmoid = 21'b111010101010110101100;
		14'b00010011001101:	sigmoid = 21'b111010101011011100100;
		14'b00010011001110:	sigmoid = 21'b111010101100000011100;
		14'b00010011001111:	sigmoid = 21'b111010101100101010100;
		14'b00010011010000:	sigmoid = 21'b111010101101010001011;
		14'b00010011010001:	sigmoid = 21'b111010101101111000001;
		14'b00010011010010:	sigmoid = 21'b111010101110011110111;
		14'b00010011010011:	sigmoid = 21'b111010101111000101100;
		14'b00010011010100:	sigmoid = 21'b111010101111101100001;
		14'b00010011010101:	sigmoid = 21'b111010110000010010110;
		14'b00010011010110:	sigmoid = 21'b111010110000111001010;
		14'b00010011010111:	sigmoid = 21'b111010110001011111101;
		14'b00010011011000:	sigmoid = 21'b111010110010000110000;
		14'b00010011011001:	sigmoid = 21'b111010110010101100011;
		14'b00010011011010:	sigmoid = 21'b111010110011010010101;
		14'b00010011011011:	sigmoid = 21'b111010110011111000110;
		14'b00010011011100:	sigmoid = 21'b111010110100011110111;
		14'b00010011011101:	sigmoid = 21'b111010110101000100111;
		14'b00010011011110:	sigmoid = 21'b111010110101101010111;
		14'b00010011011111:	sigmoid = 21'b111010110110010000111;
		14'b00010011100000:	sigmoid = 21'b111010110110110110110;
		14'b00010011100001:	sigmoid = 21'b111010110111011100100;
		14'b00010011100010:	sigmoid = 21'b111010111000000010010;
		14'b00010011100011:	sigmoid = 21'b111010111000101000000;
		14'b00010011100100:	sigmoid = 21'b111010111001001101100;
		14'b00010011100101:	sigmoid = 21'b111010111001110011001;
		14'b00010011100110:	sigmoid = 21'b111010111010011000101;
		14'b00010011100111:	sigmoid = 21'b111010111010111110000;
		14'b00010011101000:	sigmoid = 21'b111010111011100011011;
		14'b00010011101001:	sigmoid = 21'b111010111100001000110;
		14'b00010011101010:	sigmoid = 21'b111010111100101110000;
		14'b00010011101011:	sigmoid = 21'b111010111101010011001;
		14'b00010011101100:	sigmoid = 21'b111010111101111000010;
		14'b00010011101101:	sigmoid = 21'b111010111110011101011;
		14'b00010011101110:	sigmoid = 21'b111010111111000010011;
		14'b00010011101111:	sigmoid = 21'b111010111111100111011;
		14'b00010011110000:	sigmoid = 21'b111011000000001100010;
		14'b00010011110001:	sigmoid = 21'b111011000000110001000;
		14'b00010011110010:	sigmoid = 21'b111011000001010101110;
		14'b00010011110011:	sigmoid = 21'b111011000001111010100;
		14'b00010011110100:	sigmoid = 21'b111011000010011111001;
		14'b00010011110101:	sigmoid = 21'b111011000011000011110;
		14'b00010011110110:	sigmoid = 21'b111011000011101000010;
		14'b00010011110111:	sigmoid = 21'b111011000100001100110;
		14'b00010011111000:	sigmoid = 21'b111011000100110001001;
		14'b00010011111001:	sigmoid = 21'b111011000101010101100;
		14'b00010011111010:	sigmoid = 21'b111011000101111001110;
		14'b00010011111011:	sigmoid = 21'b111011000110011110000;
		14'b00010011111100:	sigmoid = 21'b111011000111000010001;
		14'b00010011111101:	sigmoid = 21'b111011000111100110010;
		14'b00010011111110:	sigmoid = 21'b111011001000001010010;
		14'b00010011111111:	sigmoid = 21'b111011001000101110010;
		14'b00010100000000:	sigmoid = 21'b111011001001010010001;
		14'b00010100000001:	sigmoid = 21'b111011001001110110000;
		14'b00010100000010:	sigmoid = 21'b111011001010011001111;
		14'b00010100000011:	sigmoid = 21'b111011001010111101101;
		14'b00010100000100:	sigmoid = 21'b111011001011100001010;
		14'b00010100000101:	sigmoid = 21'b111011001100000100111;
		14'b00010100000110:	sigmoid = 21'b111011001100101000100;
		14'b00010100000111:	sigmoid = 21'b111011001101001100000;
		14'b00010100001000:	sigmoid = 21'b111011001101101111011;
		14'b00010100001001:	sigmoid = 21'b111011001110010010110;
		14'b00010100001010:	sigmoid = 21'b111011001110110110001;
		14'b00010100001011:	sigmoid = 21'b111011001111011001011;
		14'b00010100001100:	sigmoid = 21'b111011001111111100101;
		14'b00010100001101:	sigmoid = 21'b111011010000011111110;
		14'b00010100001110:	sigmoid = 21'b111011010001000010111;
		14'b00010100001111:	sigmoid = 21'b111011010001100101111;
		14'b00010100010000:	sigmoid = 21'b111011010010001000111;
		14'b00010100010001:	sigmoid = 21'b111011010010101011111;
		14'b00010100010010:	sigmoid = 21'b111011010011001110110;
		14'b00010100010011:	sigmoid = 21'b111011010011110001100;
		14'b00010100010100:	sigmoid = 21'b111011010100010100010;
		14'b00010100010101:	sigmoid = 21'b111011010100110110111;
		14'b00010100010110:	sigmoid = 21'b111011010101011001101;
		14'b00010100010111:	sigmoid = 21'b111011010101111100001;
		14'b00010100011000:	sigmoid = 21'b111011010110011110101;
		14'b00010100011001:	sigmoid = 21'b111011010111000001001;
		14'b00010100011010:	sigmoid = 21'b111011010111100011100;
		14'b00010100011011:	sigmoid = 21'b111011011000000101111;
		14'b00010100011100:	sigmoid = 21'b111011011000101000001;
		14'b00010100011101:	sigmoid = 21'b111011011001001010011;
		14'b00010100011110:	sigmoid = 21'b111011011001101100100;
		14'b00010100011111:	sigmoid = 21'b111011011010001110101;
		14'b00010100100000:	sigmoid = 21'b111011011010110000110;
		14'b00010100100001:	sigmoid = 21'b111011011011010010110;
		14'b00010100100010:	sigmoid = 21'b111011011011110100101;
		14'b00010100100011:	sigmoid = 21'b111011011100010110101;
		14'b00010100100100:	sigmoid = 21'b111011011100111000011;
		14'b00010100100101:	sigmoid = 21'b111011011101011010001;
		14'b00010100100110:	sigmoid = 21'b111011011101111011111;
		14'b00010100100111:	sigmoid = 21'b111011011110011101100;
		14'b00010100101000:	sigmoid = 21'b111011011110111111001;
		14'b00010100101001:	sigmoid = 21'b111011011111100000110;
		14'b00010100101010:	sigmoid = 21'b111011100000000010010;
		14'b00010100101011:	sigmoid = 21'b111011100000100011101;
		14'b00010100101100:	sigmoid = 21'b111011100001000101000;
		14'b00010100101101:	sigmoid = 21'b111011100001100110011;
		14'b00010100101110:	sigmoid = 21'b111011100010000111101;
		14'b00010100101111:	sigmoid = 21'b111011100010101000111;
		14'b00010100110000:	sigmoid = 21'b111011100011001010000;
		14'b00010100110001:	sigmoid = 21'b111011100011101011001;
		14'b00010100110010:	sigmoid = 21'b111011100100001100001;
		14'b00010100110011:	sigmoid = 21'b111011100100101101001;
		14'b00010100110100:	sigmoid = 21'b111011100101001110000;
		14'b00010100110101:	sigmoid = 21'b111011100101101111000;
		14'b00010100110110:	sigmoid = 21'b111011100110001111110;
		14'b00010100110111:	sigmoid = 21'b111011100110110000100;
		14'b00010100111000:	sigmoid = 21'b111011100111010001010;
		14'b00010100111001:	sigmoid = 21'b111011100111110001111;
		14'b00010100111010:	sigmoid = 21'b111011101000010010100;
		14'b00010100111011:	sigmoid = 21'b111011101000110011000;
		14'b00010100111100:	sigmoid = 21'b111011101001010011100;
		14'b00010100111101:	sigmoid = 21'b111011101001110100000;
		14'b00010100111110:	sigmoid = 21'b111011101010010100011;
		14'b00010100111111:	sigmoid = 21'b111011101010110100110;
		14'b00010101000000:	sigmoid = 21'b111011101011010101000;
		14'b00010101000001:	sigmoid = 21'b111011101011110101010;
		14'b00010101000010:	sigmoid = 21'b111011101100010101011;
		14'b00010101000011:	sigmoid = 21'b111011101100110101100;
		14'b00010101000100:	sigmoid = 21'b111011101101010101100;
		14'b00010101000101:	sigmoid = 21'b111011101101110101100;
		14'b00010101000110:	sigmoid = 21'b111011101110010101100;
		14'b00010101000111:	sigmoid = 21'b111011101110110101011;
		14'b00010101001000:	sigmoid = 21'b111011101111010101010;
		14'b00010101001001:	sigmoid = 21'b111011101111110101000;
		14'b00010101001010:	sigmoid = 21'b111011110000010100110;
		14'b00010101001011:	sigmoid = 21'b111011110000110100011;
		14'b00010101001100:	sigmoid = 21'b111011110001010100000;
		14'b00010101001101:	sigmoid = 21'b111011110001110011101;
		14'b00010101001110:	sigmoid = 21'b111011110010010011001;
		14'b00010101001111:	sigmoid = 21'b111011110010110010101;
		14'b00010101010000:	sigmoid = 21'b111011110011010010000;
		14'b00010101010001:	sigmoid = 21'b111011110011110001011;
		14'b00010101010010:	sigmoid = 21'b111011110100010000110;
		14'b00010101010011:	sigmoid = 21'b111011110100110000000;
		14'b00010101010100:	sigmoid = 21'b111011110101001111001;
		14'b00010101010101:	sigmoid = 21'b111011110101101110010;
		14'b00010101010110:	sigmoid = 21'b111011110110001101011;
		14'b00010101010111:	sigmoid = 21'b111011110110101100011;
		14'b00010101011000:	sigmoid = 21'b111011110111001011011;
		14'b00010101011001:	sigmoid = 21'b111011110111101010011;
		14'b00010101011010:	sigmoid = 21'b111011111000001001010;
		14'b00010101011011:	sigmoid = 21'b111011111000101000001;
		14'b00010101011100:	sigmoid = 21'b111011111001000110111;
		14'b00010101011101:	sigmoid = 21'b111011111001100101101;
		14'b00010101011110:	sigmoid = 21'b111011111010000100010;
		14'b00010101011111:	sigmoid = 21'b111011111010100010111;
		14'b00010101100000:	sigmoid = 21'b111011111011000001011;
		14'b00010101100001:	sigmoid = 21'b111011111011100000000;
		14'b00010101100010:	sigmoid = 21'b111011111011111110011;
		14'b00010101100011:	sigmoid = 21'b111011111100011100111;
		14'b00010101100100:	sigmoid = 21'b111011111100111011010;
		14'b00010101100101:	sigmoid = 21'b111011111101011001100;
		14'b00010101100110:	sigmoid = 21'b111011111101110111110;
		14'b00010101100111:	sigmoid = 21'b111011111110010110000;
		14'b00010101101000:	sigmoid = 21'b111011111110110100001;
		14'b00010101101001:	sigmoid = 21'b111011111111010010010;
		14'b00010101101010:	sigmoid = 21'b111011111111110000010;
		14'b00010101101011:	sigmoid = 21'b111100000000001110010;
		14'b00010101101100:	sigmoid = 21'b111100000000101100010;
		14'b00010101101101:	sigmoid = 21'b111100000001001010001;
		14'b00010101101110:	sigmoid = 21'b111100000001101000000;
		14'b00010101101111:	sigmoid = 21'b111100000010000101110;
		14'b00010101110000:	sigmoid = 21'b111100000010100011100;
		14'b00010101110001:	sigmoid = 21'b111100000011000001010;
		14'b00010101110010:	sigmoid = 21'b111100000011011110111;
		14'b00010101110011:	sigmoid = 21'b111100000011111100100;
		14'b00010101110100:	sigmoid = 21'b111100000100011010000;
		14'b00010101110101:	sigmoid = 21'b111100000100110111100;
		14'b00010101110110:	sigmoid = 21'b111100000101010100111;
		14'b00010101110111:	sigmoid = 21'b111100000101110010011;
		14'b00010101111000:	sigmoid = 21'b111100000110001111101;
		14'b00010101111001:	sigmoid = 21'b111100000110101101000;
		14'b00010101111010:	sigmoid = 21'b111100000111001010010;
		14'b00010101111011:	sigmoid = 21'b111100000111100111011;
		14'b00010101111100:	sigmoid = 21'b111100001000000100100;
		14'b00010101111101:	sigmoid = 21'b111100001000100001101;
		14'b00010101111110:	sigmoid = 21'b111100001000111110101;
		14'b00010101111111:	sigmoid = 21'b111100001001011011101;
		14'b00010110000000:	sigmoid = 21'b111100001001111000101;
		14'b00010110000001:	sigmoid = 21'b111100001010010101100;
		14'b00010110000010:	sigmoid = 21'b111100001010110010011;
		14'b00010110000011:	sigmoid = 21'b111100001011001111001;
		14'b00010110000100:	sigmoid = 21'b111100001011101011111;
		14'b00010110000101:	sigmoid = 21'b111100001100001000100;
		14'b00010110000110:	sigmoid = 21'b111100001100100101001;
		14'b00010110000111:	sigmoid = 21'b111100001101000001110;
		14'b00010110001000:	sigmoid = 21'b111100001101011110011;
		14'b00010110001001:	sigmoid = 21'b111100001101111010111;
		14'b00010110001010:	sigmoid = 21'b111100001110010111010;
		14'b00010110001011:	sigmoid = 21'b111100001110110011101;
		14'b00010110001100:	sigmoid = 21'b111100001111010000000;
		14'b00010110001101:	sigmoid = 21'b111100001111101100011;
		14'b00010110001110:	sigmoid = 21'b111100010000001000101;
		14'b00010110001111:	sigmoid = 21'b111100010000100100110;
		14'b00010110010000:	sigmoid = 21'b111100010001000000111;
		14'b00010110010001:	sigmoid = 21'b111100010001011101000;
		14'b00010110010010:	sigmoid = 21'b111100010001111001001;
		14'b00010110010011:	sigmoid = 21'b111100010010010101001;
		14'b00010110010100:	sigmoid = 21'b111100010010110001000;
		14'b00010110010101:	sigmoid = 21'b111100010011001101000;
		14'b00010110010110:	sigmoid = 21'b111100010011101000111;
		14'b00010110010111:	sigmoid = 21'b111100010100000100101;
		14'b00010110011000:	sigmoid = 21'b111100010100100000011;
		14'b00010110011001:	sigmoid = 21'b111100010100111100001;
		14'b00010110011010:	sigmoid = 21'b111100010101010111110;
		14'b00010110011011:	sigmoid = 21'b111100010101110011011;
		14'b00010110011100:	sigmoid = 21'b111100010110001111000;
		14'b00010110011101:	sigmoid = 21'b111100010110101010100;
		14'b00010110011110:	sigmoid = 21'b111100010111000110000;
		14'b00010110011111:	sigmoid = 21'b111100010111100001100;
		14'b00010110100000:	sigmoid = 21'b111100010111111100111;
		14'b00010110100001:	sigmoid = 21'b111100011000011000001;
		14'b00010110100010:	sigmoid = 21'b111100011000110011100;
		14'b00010110100011:	sigmoid = 21'b111100011001001110110;
		14'b00010110100100:	sigmoid = 21'b111100011001101001111;
		14'b00010110100101:	sigmoid = 21'b111100011010000101001;
		14'b00010110100110:	sigmoid = 21'b111100011010100000001;
		14'b00010110100111:	sigmoid = 21'b111100011010111011010;
		14'b00010110101000:	sigmoid = 21'b111100011011010110010;
		14'b00010110101001:	sigmoid = 21'b111100011011110001010;
		14'b00010110101010:	sigmoid = 21'b111100011100001100001;
		14'b00010110101011:	sigmoid = 21'b111100011100100111000;
		14'b00010110101100:	sigmoid = 21'b111100011101000001110;
		14'b00010110101101:	sigmoid = 21'b111100011101011100101;
		14'b00010110101110:	sigmoid = 21'b111100011101110111010;
		14'b00010110101111:	sigmoid = 21'b111100011110010010000;
		14'b00010110110000:	sigmoid = 21'b111100011110101100101;
		14'b00010110110001:	sigmoid = 21'b111100011111000111010;
		14'b00010110110010:	sigmoid = 21'b111100011111100001110;
		14'b00010110110011:	sigmoid = 21'b111100011111111100010;
		14'b00010110110100:	sigmoid = 21'b111100100000010110110;
		14'b00010110110101:	sigmoid = 21'b111100100000110001001;
		14'b00010110110110:	sigmoid = 21'b111100100001001011100;
		14'b00010110110111:	sigmoid = 21'b111100100001100101110;
		14'b00010110111000:	sigmoid = 21'b111100100010000000001;
		14'b00010110111001:	sigmoid = 21'b111100100010011010010;
		14'b00010110111010:	sigmoid = 21'b111100100010110100100;
		14'b00010110111011:	sigmoid = 21'b111100100011001110101;
		14'b00010110111100:	sigmoid = 21'b111100100011101000101;
		14'b00010110111101:	sigmoid = 21'b111100100100000010110;
		14'b00010110111110:	sigmoid = 21'b111100100100011100110;
		14'b00010110111111:	sigmoid = 21'b111100100100110110101;
		14'b00010111000000:	sigmoid = 21'b111100100101010000101;
		14'b00010111000001:	sigmoid = 21'b111100100101101010011;
		14'b00010111000010:	sigmoid = 21'b111100100110000100010;
		14'b00010111000011:	sigmoid = 21'b111100100110011110000;
		14'b00010111000100:	sigmoid = 21'b111100100110110111110;
		14'b00010111000101:	sigmoid = 21'b111100100111010001011;
		14'b00010111000110:	sigmoid = 21'b111100100111101011000;
		14'b00010111000111:	sigmoid = 21'b111100101000000100101;
		14'b00010111001000:	sigmoid = 21'b111100101000011110010;
		14'b00010111001001:	sigmoid = 21'b111100101000110111110;
		14'b00010111001010:	sigmoid = 21'b111100101001010001001;
		14'b00010111001011:	sigmoid = 21'b111100101001101010101;
		14'b00010111001100:	sigmoid = 21'b111100101010000011111;
		14'b00010111001101:	sigmoid = 21'b111100101010011101010;
		14'b00010111001110:	sigmoid = 21'b111100101010110110100;
		14'b00010111001111:	sigmoid = 21'b111100101011001111110;
		14'b00010111010000:	sigmoid = 21'b111100101011101001000;
		14'b00010111010001:	sigmoid = 21'b111100101100000010001;
		14'b00010111010010:	sigmoid = 21'b111100101100011011010;
		14'b00010111010011:	sigmoid = 21'b111100101100110100010;
		14'b00010111010100:	sigmoid = 21'b111100101101001101010;
		14'b00010111010101:	sigmoid = 21'b111100101101100110010;
		14'b00010111010110:	sigmoid = 21'b111100101101111111001;
		14'b00010111010111:	sigmoid = 21'b111100101110011000001;
		14'b00010111011000:	sigmoid = 21'b111100101110110000111;
		14'b00010111011001:	sigmoid = 21'b111100101111001001110;
		14'b00010111011010:	sigmoid = 21'b111100101111100010100;
		14'b00010111011011:	sigmoid = 21'b111100101111111011001;
		14'b00010111011100:	sigmoid = 21'b111100110000010011111;
		14'b00010111011101:	sigmoid = 21'b111100110000101100100;
		14'b00010111011110:	sigmoid = 21'b111100110001000101000;
		14'b00010111011111:	sigmoid = 21'b111100110001011101101;
		14'b00010111100000:	sigmoid = 21'b111100110001110110001;
		14'b00010111100001:	sigmoid = 21'b111100110010001110100;
		14'b00010111100010:	sigmoid = 21'b111100110010100110111;
		14'b00010111100011:	sigmoid = 21'b111100110010111111010;
		14'b00010111100100:	sigmoid = 21'b111100110011010111101;
		14'b00010111100101:	sigmoid = 21'b111100110011101111111;
		14'b00010111100110:	sigmoid = 21'b111100110100001000001;
		14'b00010111100111:	sigmoid = 21'b111100110100100000011;
		14'b00010111101000:	sigmoid = 21'b111100110100111000100;
		14'b00010111101001:	sigmoid = 21'b111100110101010000101;
		14'b00010111101010:	sigmoid = 21'b111100110101101000101;
		14'b00010111101011:	sigmoid = 21'b111100110110000000101;
		14'b00010111101100:	sigmoid = 21'b111100110110011000101;
		14'b00010111101101:	sigmoid = 21'b111100110110110000101;
		14'b00010111101110:	sigmoid = 21'b111100110111001000100;
		14'b00010111101111:	sigmoid = 21'b111100110111100000011;
		14'b00010111110000:	sigmoid = 21'b111100110111111000001;
		14'b00010111110001:	sigmoid = 21'b111100111000001111111;
		14'b00010111110010:	sigmoid = 21'b111100111000100111101;
		14'b00010111110011:	sigmoid = 21'b111100111000111111011;
		14'b00010111110100:	sigmoid = 21'b111100111001010111000;
		14'b00010111110101:	sigmoid = 21'b111100111001101110101;
		14'b00010111110110:	sigmoid = 21'b111100111010000110001;
		14'b00010111110111:	sigmoid = 21'b111100111010011101110;
		14'b00010111111000:	sigmoid = 21'b111100111010110101001;
		14'b00010111111001:	sigmoid = 21'b111100111011001100101;
		14'b00010111111010:	sigmoid = 21'b111100111011100100000;
		14'b00010111111011:	sigmoid = 21'b111100111011111011011;
		14'b00010111111100:	sigmoid = 21'b111100111100010010101;
		14'b00010111111101:	sigmoid = 21'b111100111100101010000;
		14'b00010111111110:	sigmoid = 21'b111100111101000001001;
		14'b00010111111111:	sigmoid = 21'b111100111101011000011;
		14'b00011000000000:	sigmoid = 21'b111100111101101111100;
		14'b00011000000001:	sigmoid = 21'b111100111110000110101;
		14'b00011000000010:	sigmoid = 21'b111100111110011101110;
		14'b00011000000011:	sigmoid = 21'b111100111110110100110;
		14'b00011000000100:	sigmoid = 21'b111100111111001011110;
		14'b00011000000101:	sigmoid = 21'b111100111111100010101;
		14'b00011000000110:	sigmoid = 21'b111100111111111001101;
		14'b00011000000111:	sigmoid = 21'b111101000000010000100;
		14'b00011000001000:	sigmoid = 21'b111101000000100111010;
		14'b00011000001001:	sigmoid = 21'b111101000000111110000;
		14'b00011000001010:	sigmoid = 21'b111101000001010100110;
		14'b00011000001011:	sigmoid = 21'b111101000001101011100;
		14'b00011000001100:	sigmoid = 21'b111101000010000010001;
		14'b00011000001101:	sigmoid = 21'b111101000010011000110;
		14'b00011000001110:	sigmoid = 21'b111101000010101111011;
		14'b00011000001111:	sigmoid = 21'b111101000011000101111;
		14'b00011000010000:	sigmoid = 21'b111101000011011100011;
		14'b00011000010001:	sigmoid = 21'b111101000011110010111;
		14'b00011000010010:	sigmoid = 21'b111101000100001001011;
		14'b00011000010011:	sigmoid = 21'b111101000100011111110;
		14'b00011000010100:	sigmoid = 21'b111101000100110110000;
		14'b00011000010101:	sigmoid = 21'b111101000101001100011;
		14'b00011000010110:	sigmoid = 21'b111101000101100010101;
		14'b00011000010111:	sigmoid = 21'b111101000101111000111;
		14'b00011000011000:	sigmoid = 21'b111101000110001111000;
		14'b00011000011001:	sigmoid = 21'b111101000110100101001;
		14'b00011000011010:	sigmoid = 21'b111101000110111011010;
		14'b00011000011011:	sigmoid = 21'b111101000111010001011;
		14'b00011000011100:	sigmoid = 21'b111101000111100111011;
		14'b00011000011101:	sigmoid = 21'b111101000111111101011;
		14'b00011000011110:	sigmoid = 21'b111101001000010011011;
		14'b00011000011111:	sigmoid = 21'b111101001000101001010;
		14'b00011000100000:	sigmoid = 21'b111101001000111111001;
		14'b00011000100001:	sigmoid = 21'b111101001001010101000;
		14'b00011000100010:	sigmoid = 21'b111101001001101010110;
		14'b00011000100011:	sigmoid = 21'b111101001010000000100;
		14'b00011000100100:	sigmoid = 21'b111101001010010110010;
		14'b00011000100101:	sigmoid = 21'b111101001010101011111;
		14'b00011000100110:	sigmoid = 21'b111101001011000001100;
		14'b00011000100111:	sigmoid = 21'b111101001011010111001;
		14'b00011000101000:	sigmoid = 21'b111101001011101100110;
		14'b00011000101001:	sigmoid = 21'b111101001100000010010;
		14'b00011000101010:	sigmoid = 21'b111101001100010111110;
		14'b00011000101011:	sigmoid = 21'b111101001100101101001;
		14'b00011000101100:	sigmoid = 21'b111101001101000010101;
		14'b00011000101101:	sigmoid = 21'b111101001101011000000;
		14'b00011000101110:	sigmoid = 21'b111101001101101101010;
		14'b00011000101111:	sigmoid = 21'b111101001110000010101;
		14'b00011000110000:	sigmoid = 21'b111101001110010111111;
		14'b00011000110001:	sigmoid = 21'b111101001110101101001;
		14'b00011000110010:	sigmoid = 21'b111101001111000010010;
		14'b00011000110011:	sigmoid = 21'b111101001111010111011;
		14'b00011000110100:	sigmoid = 21'b111101001111101100100;
		14'b00011000110101:	sigmoid = 21'b111101010000000001101;
		14'b00011000110110:	sigmoid = 21'b111101010000010110101;
		14'b00011000110111:	sigmoid = 21'b111101010000101011101;
		14'b00011000111000:	sigmoid = 21'b111101010001000000101;
		14'b00011000111001:	sigmoid = 21'b111101010001010101100;
		14'b00011000111010:	sigmoid = 21'b111101010001101010011;
		14'b00011000111011:	sigmoid = 21'b111101010001111111010;
		14'b00011000111100:	sigmoid = 21'b111101010010010100000;
		14'b00011000111101:	sigmoid = 21'b111101010010101000110;
		14'b00011000111110:	sigmoid = 21'b111101010010111101100;
		14'b00011000111111:	sigmoid = 21'b111101010011010010010;
		14'b00011001000000:	sigmoid = 21'b111101010011100110111;
		14'b00011001000001:	sigmoid = 21'b111101010011111011100;
		14'b00011001000010:	sigmoid = 21'b111101010100010000001;
		14'b00011001000011:	sigmoid = 21'b111101010100100100101;
		14'b00011001000100:	sigmoid = 21'b111101010100111001001;
		14'b00011001000101:	sigmoid = 21'b111101010101001101101;
		14'b00011001000110:	sigmoid = 21'b111101010101100010001;
		14'b00011001000111:	sigmoid = 21'b111101010101110110100;
		14'b00011001001000:	sigmoid = 21'b111101010110001010111;
		14'b00011001001001:	sigmoid = 21'b111101010110011111001;
		14'b00011001001010:	sigmoid = 21'b111101010110110011100;
		14'b00011001001011:	sigmoid = 21'b111101010111000111110;
		14'b00011001001100:	sigmoid = 21'b111101010111011100000;
		14'b00011001001101:	sigmoid = 21'b111101010111110000001;
		14'b00011001001110:	sigmoid = 21'b111101011000000100010;
		14'b00011001001111:	sigmoid = 21'b111101011000011000011;
		14'b00011001010000:	sigmoid = 21'b111101011000101100100;
		14'b00011001010001:	sigmoid = 21'b111101011001000000100;
		14'b00011001010010:	sigmoid = 21'b111101011001010100100;
		14'b00011001010011:	sigmoid = 21'b111101011001101000100;
		14'b00011001010100:	sigmoid = 21'b111101011001111100011;
		14'b00011001010101:	sigmoid = 21'b111101011010010000011;
		14'b00011001010110:	sigmoid = 21'b111101011010100100001;
		14'b00011001010111:	sigmoid = 21'b111101011010111000000;
		14'b00011001011000:	sigmoid = 21'b111101011011001011110;
		14'b00011001011001:	sigmoid = 21'b111101011011011111100;
		14'b00011001011010:	sigmoid = 21'b111101011011110011010;
		14'b00011001011011:	sigmoid = 21'b111101011100000111000;
		14'b00011001011100:	sigmoid = 21'b111101011100011010101;
		14'b00011001011101:	sigmoid = 21'b111101011100101110010;
		14'b00011001011110:	sigmoid = 21'b111101011101000001110;
		14'b00011001011111:	sigmoid = 21'b111101011101010101011;
		14'b00011001100000:	sigmoid = 21'b111101011101101000111;
		14'b00011001100001:	sigmoid = 21'b111101011101111100011;
		14'b00011001100010:	sigmoid = 21'b111101011110001111110;
		14'b00011001100011:	sigmoid = 21'b111101011110100011001;
		14'b00011001100100:	sigmoid = 21'b111101011110110110100;
		14'b00011001100101:	sigmoid = 21'b111101011111001001111;
		14'b00011001100110:	sigmoid = 21'b111101011111011101001;
		14'b00011001100111:	sigmoid = 21'b111101011111110000011;
		14'b00011001101000:	sigmoid = 21'b111101100000000011101;
		14'b00011001101001:	sigmoid = 21'b111101100000010110111;
		14'b00011001101010:	sigmoid = 21'b111101100000101010000;
		14'b00011001101011:	sigmoid = 21'b111101100000111101001;
		14'b00011001101100:	sigmoid = 21'b111101100001010000010;
		14'b00011001101101:	sigmoid = 21'b111101100001100011010;
		14'b00011001101110:	sigmoid = 21'b111101100001110110011;
		14'b00011001101111:	sigmoid = 21'b111101100010001001010;
		14'b00011001110000:	sigmoid = 21'b111101100010011100010;
		14'b00011001110001:	sigmoid = 21'b111101100010101111001;
		14'b00011001110010:	sigmoid = 21'b111101100011000010000;
		14'b00011001110011:	sigmoid = 21'b111101100011010100111;
		14'b00011001110100:	sigmoid = 21'b111101100011100111110;
		14'b00011001110101:	sigmoid = 21'b111101100011111010100;
		14'b00011001110110:	sigmoid = 21'b111101100100001101010;
		14'b00011001110111:	sigmoid = 21'b111101100100100000000;
		14'b00011001111000:	sigmoid = 21'b111101100100110010101;
		14'b00011001111001:	sigmoid = 21'b111101100101000101011;
		14'b00011001111010:	sigmoid = 21'b111101100101010111111;
		14'b00011001111011:	sigmoid = 21'b111101100101101010100;
		14'b00011001111100:	sigmoid = 21'b111101100101111101000;
		14'b00011001111101:	sigmoid = 21'b111101100110001111101;
		14'b00011001111110:	sigmoid = 21'b111101100110100010000;
		14'b00011001111111:	sigmoid = 21'b111101100110110100100;
		14'b00011010000000:	sigmoid = 21'b111101100111000110111;
		14'b00011010000001:	sigmoid = 21'b111101100111011001010;
		14'b00011010000010:	sigmoid = 21'b111101100111101011101;
		14'b00011010000011:	sigmoid = 21'b111101100111111110000;
		14'b00011010000100:	sigmoid = 21'b111101101000010000010;
		14'b00011010000101:	sigmoid = 21'b111101101000100010100;
		14'b00011010000110:	sigmoid = 21'b111101101000110100110;
		14'b00011010000111:	sigmoid = 21'b111101101001000110111;
		14'b00011010001000:	sigmoid = 21'b111101101001011001000;
		14'b00011010001001:	sigmoid = 21'b111101101001101011001;
		14'b00011010001010:	sigmoid = 21'b111101101001111101010;
		14'b00011010001011:	sigmoid = 21'b111101101010001111010;
		14'b00011010001100:	sigmoid = 21'b111101101010100001011;
		14'b00011010001101:	sigmoid = 21'b111101101010110011010;
		14'b00011010001110:	sigmoid = 21'b111101101011000101010;
		14'b00011010001111:	sigmoid = 21'b111101101011010111001;
		14'b00011010010000:	sigmoid = 21'b111101101011101001001;
		14'b00011010010001:	sigmoid = 21'b111101101011111010111;
		14'b00011010010010:	sigmoid = 21'b111101101100001100110;
		14'b00011010010011:	sigmoid = 21'b111101101100011110100;
		14'b00011010010100:	sigmoid = 21'b111101101100110000010;
		14'b00011010010101:	sigmoid = 21'b111101101101000010000;
		14'b00011010010110:	sigmoid = 21'b111101101101010011110;
		14'b00011010010111:	sigmoid = 21'b111101101101100101011;
		14'b00011010011000:	sigmoid = 21'b111101101101110111000;
		14'b00011010011001:	sigmoid = 21'b111101101110001000101;
		14'b00011010011010:	sigmoid = 21'b111101101110011010001;
		14'b00011010011011:	sigmoid = 21'b111101101110101011110;
		14'b00011010011100:	sigmoid = 21'b111101101110111101010;
		14'b00011010011101:	sigmoid = 21'b111101101111001110110;
		14'b00011010011110:	sigmoid = 21'b111101101111100000001;
		14'b00011010011111:	sigmoid = 21'b111101101111110001100;
		14'b00011010100000:	sigmoid = 21'b111101110000000010111;
		14'b00011010100001:	sigmoid = 21'b111101110000010100010;
		14'b00011010100010:	sigmoid = 21'b111101110000100101101;
		14'b00011010100011:	sigmoid = 21'b111101110000110110111;
		14'b00011010100100:	sigmoid = 21'b111101110001001000001;
		14'b00011010100101:	sigmoid = 21'b111101110001011001011;
		14'b00011010100110:	sigmoid = 21'b111101110001101010100;
		14'b00011010100111:	sigmoid = 21'b111101110001111011110;
		14'b00011010101000:	sigmoid = 21'b111101110010001100111;
		14'b00011010101001:	sigmoid = 21'b111101110010011101111;
		14'b00011010101010:	sigmoid = 21'b111101110010101111000;
		14'b00011010101011:	sigmoid = 21'b111101110011000000000;
		14'b00011010101100:	sigmoid = 21'b111101110011010001000;
		14'b00011010101101:	sigmoid = 21'b111101110011100010000;
		14'b00011010101110:	sigmoid = 21'b111101110011110010111;
		14'b00011010101111:	sigmoid = 21'b111101110100000011111;
		14'b00011010110000:	sigmoid = 21'b111101110100010100110;
		14'b00011010110001:	sigmoid = 21'b111101110100100101101;
		14'b00011010110010:	sigmoid = 21'b111101110100110110011;
		14'b00011010110011:	sigmoid = 21'b111101110101000111001;
		14'b00011010110100:	sigmoid = 21'b111101110101010111111;
		14'b00011010110101:	sigmoid = 21'b111101110101101000101;
		14'b00011010110110:	sigmoid = 21'b111101110101111001011;
		14'b00011010110111:	sigmoid = 21'b111101110110001010000;
		14'b00011010111000:	sigmoid = 21'b111101110110011010101;
		14'b00011010111001:	sigmoid = 21'b111101110110101011010;
		14'b00011010111010:	sigmoid = 21'b111101110110111011111;
		14'b00011010111011:	sigmoid = 21'b111101110111001100011;
		14'b00011010111100:	sigmoid = 21'b111101110111011100111;
		14'b00011010111101:	sigmoid = 21'b111101110111101101011;
		14'b00011010111110:	sigmoid = 21'b111101110111111101111;
		14'b00011010111111:	sigmoid = 21'b111101111000001110010;
		14'b00011011000000:	sigmoid = 21'b111101111000011110101;
		14'b00011011000001:	sigmoid = 21'b111101111000101111000;
		14'b00011011000010:	sigmoid = 21'b111101111000111111011;
		14'b00011011000011:	sigmoid = 21'b111101111001001111101;
		14'b00011011000100:	sigmoid = 21'b111101111001011111111;
		14'b00011011000101:	sigmoid = 21'b111101111001110000001;
		14'b00011011000110:	sigmoid = 21'b111101111010000000011;
		14'b00011011000111:	sigmoid = 21'b111101111010010000101;
		14'b00011011001000:	sigmoid = 21'b111101111010100000110;
		14'b00011011001001:	sigmoid = 21'b111101111010110000111;
		14'b00011011001010:	sigmoid = 21'b111101111011000001000;
		14'b00011011001011:	sigmoid = 21'b111101111011010001000;
		14'b00011011001100:	sigmoid = 21'b111101111011100001001;
		14'b00011011001101:	sigmoid = 21'b111101111011110001001;
		14'b00011011001110:	sigmoid = 21'b111101111100000001000;
		14'b00011011001111:	sigmoid = 21'b111101111100010001000;
		14'b00011011010000:	sigmoid = 21'b111101111100100000111;
		14'b00011011010001:	sigmoid = 21'b111101111100110000111;
		14'b00011011010010:	sigmoid = 21'b111101111101000000110;
		14'b00011011010011:	sigmoid = 21'b111101111101010000100;
		14'b00011011010100:	sigmoid = 21'b111101111101100000011;
		14'b00011011010101:	sigmoid = 21'b111101111101110000001;
		14'b00011011010110:	sigmoid = 21'b111101111101111111111;
		14'b00011011010111:	sigmoid = 21'b111101111110001111101;
		14'b00011011011000:	sigmoid = 21'b111101111110011111010;
		14'b00011011011001:	sigmoid = 21'b111101111110101110111;
		14'b00011011011010:	sigmoid = 21'b111101111110111110101;
		14'b00011011011011:	sigmoid = 21'b111101111111001110001;
		14'b00011011011100:	sigmoid = 21'b111101111111011101110;
		14'b00011011011101:	sigmoid = 21'b111101111111101101010;
		14'b00011011011110:	sigmoid = 21'b111101111111111100111;
		14'b00011011011111:	sigmoid = 21'b111110000000001100010;
		14'b00011011100000:	sigmoid = 21'b111110000000011011110;
		14'b00011011100001:	sigmoid = 21'b111110000000101011010;
		14'b00011011100010:	sigmoid = 21'b111110000000111010101;
		14'b00011011100011:	sigmoid = 21'b111110000001001010000;
		14'b00011011100100:	sigmoid = 21'b111110000001011001011;
		14'b00011011100101:	sigmoid = 21'b111110000001101000101;
		14'b00011011100110:	sigmoid = 21'b111110000001111000000;
		14'b00011011100111:	sigmoid = 21'b111110000010000111010;
		14'b00011011101000:	sigmoid = 21'b111110000010010110100;
		14'b00011011101001:	sigmoid = 21'b111110000010100101101;
		14'b00011011101010:	sigmoid = 21'b111110000010110100111;
		14'b00011011101011:	sigmoid = 21'b111110000011000100000;
		14'b00011011101100:	sigmoid = 21'b111110000011010011001;
		14'b00011011101101:	sigmoid = 21'b111110000011100010010;
		14'b00011011101110:	sigmoid = 21'b111110000011110001010;
		14'b00011011101111:	sigmoid = 21'b111110000100000000011;
		14'b00011011110000:	sigmoid = 21'b111110000100001111011;
		14'b00011011110001:	sigmoid = 21'b111110000100011110011;
		14'b00011011110010:	sigmoid = 21'b111110000100101101011;
		14'b00011011110011:	sigmoid = 21'b111110000100111100010;
		14'b00011011110100:	sigmoid = 21'b111110000101001011001;
		14'b00011011110101:	sigmoid = 21'b111110000101011010000;
		14'b00011011110110:	sigmoid = 21'b111110000101101000111;
		14'b00011011110111:	sigmoid = 21'b111110000101110111110;
		14'b00011011111000:	sigmoid = 21'b111110000110000110100;
		14'b00011011111001:	sigmoid = 21'b111110000110010101010;
		14'b00011011111010:	sigmoid = 21'b111110000110100100000;
		14'b00011011111011:	sigmoid = 21'b111110000110110010110;
		14'b00011011111100:	sigmoid = 21'b111110000111000001011;
		14'b00011011111101:	sigmoid = 21'b111110000111010000001;
		14'b00011011111110:	sigmoid = 21'b111110000111011110110;
		14'b00011011111111:	sigmoid = 21'b111110000111101101011;
		14'b00011100000000:	sigmoid = 21'b111110000111111011111;
		14'b00011100000001:	sigmoid = 21'b111110001000001010100;
		14'b00011100000010:	sigmoid = 21'b111110001000011001000;
		14'b00011100000011:	sigmoid = 21'b111110001000100111100;
		14'b00011100000100:	sigmoid = 21'b111110001000110110000;
		14'b00011100000101:	sigmoid = 21'b111110001001000100011;
		14'b00011100000110:	sigmoid = 21'b111110001001010010111;
		14'b00011100000111:	sigmoid = 21'b111110001001100001010;
		14'b00011100001000:	sigmoid = 21'b111110001001101111101;
		14'b00011100001001:	sigmoid = 21'b111110001001111110000;
		14'b00011100001010:	sigmoid = 21'b111110001010001100010;
		14'b00011100001011:	sigmoid = 21'b111110001010011010100;
		14'b00011100001100:	sigmoid = 21'b111110001010101000110;
		14'b00011100001101:	sigmoid = 21'b111110001010110111000;
		14'b00011100001110:	sigmoid = 21'b111110001011000101010;
		14'b00011100001111:	sigmoid = 21'b111110001011010011100;
		14'b00011100010000:	sigmoid = 21'b111110001011100001101;
		14'b00011100010001:	sigmoid = 21'b111110001011101111110;
		14'b00011100010010:	sigmoid = 21'b111110001011111101111;
		14'b00011100010011:	sigmoid = 21'b111110001100001011111;
		14'b00011100010100:	sigmoid = 21'b111110001100011010000;
		14'b00011100010101:	sigmoid = 21'b111110001100101000000;
		14'b00011100010110:	sigmoid = 21'b111110001100110110000;
		14'b00011100010111:	sigmoid = 21'b111110001101000100000;
		14'b00011100011000:	sigmoid = 21'b111110001101010001111;
		14'b00011100011001:	sigmoid = 21'b111110001101011111111;
		14'b00011100011010:	sigmoid = 21'b111110001101101101110;
		14'b00011100011011:	sigmoid = 21'b111110001101111011101;
		14'b00011100011100:	sigmoid = 21'b111110001110001001100;
		14'b00011100011101:	sigmoid = 21'b111110001110010111010;
		14'b00011100011110:	sigmoid = 21'b111110001110100101001;
		14'b00011100011111:	sigmoid = 21'b111110001110110010111;
		14'b00011100100000:	sigmoid = 21'b111110001111000000101;
		14'b00011100100001:	sigmoid = 21'b111110001111001110011;
		14'b00011100100010:	sigmoid = 21'b111110001111011100000;
		14'b00011100100011:	sigmoid = 21'b111110001111101001110;
		14'b00011100100100:	sigmoid = 21'b111110001111110111011;
		14'b00011100100101:	sigmoid = 21'b111110010000000101000;
		14'b00011100100110:	sigmoid = 21'b111110010000010010101;
		14'b00011100100111:	sigmoid = 21'b111110010000100000001;
		14'b00011100101000:	sigmoid = 21'b111110010000101101101;
		14'b00011100101001:	sigmoid = 21'b111110010000111011010;
		14'b00011100101010:	sigmoid = 21'b111110010001001000110;
		14'b00011100101011:	sigmoid = 21'b111110010001010110001;
		14'b00011100101100:	sigmoid = 21'b111110010001100011101;
		14'b00011100101101:	sigmoid = 21'b111110010001110001000;
		14'b00011100101110:	sigmoid = 21'b111110010001111110011;
		14'b00011100101111:	sigmoid = 21'b111110010010001011110;
		14'b00011100110000:	sigmoid = 21'b111110010010011001001;
		14'b00011100110001:	sigmoid = 21'b111110010010100110100;
		14'b00011100110010:	sigmoid = 21'b111110010010110011110;
		14'b00011100110011:	sigmoid = 21'b111110010011000001000;
		14'b00011100110100:	sigmoid = 21'b111110010011001110010;
		14'b00011100110101:	sigmoid = 21'b111110010011011011100;
		14'b00011100110110:	sigmoid = 21'b111110010011101000110;
		14'b00011100110111:	sigmoid = 21'b111110010011110101111;
		14'b00011100111000:	sigmoid = 21'b111110010100000011000;
		14'b00011100111001:	sigmoid = 21'b111110010100010000001;
		14'b00011100111010:	sigmoid = 21'b111110010100011101010;
		14'b00011100111011:	sigmoid = 21'b111110010100101010011;
		14'b00011100111100:	sigmoid = 21'b111110010100110111011;
		14'b00011100111101:	sigmoid = 21'b111110010101000100011;
		14'b00011100111110:	sigmoid = 21'b111110010101010001011;
		14'b00011100111111:	sigmoid = 21'b111110010101011110011;
		14'b00011101000000:	sigmoid = 21'b111110010101101011011;
		14'b00011101000001:	sigmoid = 21'b111110010101111000010;
		14'b00011101000010:	sigmoid = 21'b111110010110000101010;
		14'b00011101000011:	sigmoid = 21'b111110010110010010001;
		14'b00011101000100:	sigmoid = 21'b111110010110011111000;
		14'b00011101000101:	sigmoid = 21'b111110010110101011110;
		14'b00011101000110:	sigmoid = 21'b111110010110111000101;
		14'b00011101000111:	sigmoid = 21'b111110010111000101011;
		14'b00011101001000:	sigmoid = 21'b111110010111010010001;
		14'b00011101001001:	sigmoid = 21'b111110010111011110111;
		14'b00011101001010:	sigmoid = 21'b111110010111101011101;
		14'b00011101001011:	sigmoid = 21'b111110010111111000011;
		14'b00011101001100:	sigmoid = 21'b111110011000000101000;
		14'b00011101001101:	sigmoid = 21'b111110011000010001101;
		14'b00011101001110:	sigmoid = 21'b111110011000011110010;
		14'b00011101001111:	sigmoid = 21'b111110011000101010111;
		14'b00011101010000:	sigmoid = 21'b111110011000110111100;
		14'b00011101010001:	sigmoid = 21'b111110011001000100000;
		14'b00011101010010:	sigmoid = 21'b111110011001010000100;
		14'b00011101010011:	sigmoid = 21'b111110011001011101000;
		14'b00011101010100:	sigmoid = 21'b111110011001101001100;
		14'b00011101010101:	sigmoid = 21'b111110011001110110000;
		14'b00011101010110:	sigmoid = 21'b111110011010000010100;
		14'b00011101010111:	sigmoid = 21'b111110011010001110111;
		14'b00011101011000:	sigmoid = 21'b111110011010011011010;
		14'b00011101011001:	sigmoid = 21'b111110011010100111101;
		14'b00011101011010:	sigmoid = 21'b111110011010110100000;
		14'b00011101011011:	sigmoid = 21'b111110011011000000010;
		14'b00011101011100:	sigmoid = 21'b111110011011001100101;
		14'b00011101011101:	sigmoid = 21'b111110011011011000111;
		14'b00011101011110:	sigmoid = 21'b111110011011100101001;
		14'b00011101011111:	sigmoid = 21'b111110011011110001011;
		14'b00011101100000:	sigmoid = 21'b111110011011111101101;
		14'b00011101100001:	sigmoid = 21'b111110011100001001110;
		14'b00011101100010:	sigmoid = 21'b111110011100010101111;
		14'b00011101100011:	sigmoid = 21'b111110011100100010001;
		14'b00011101100100:	sigmoid = 21'b111110011100101110001;
		14'b00011101100101:	sigmoid = 21'b111110011100111010010;
		14'b00011101100110:	sigmoid = 21'b111110011101000110011;
		14'b00011101100111:	sigmoid = 21'b111110011101010010011;
		14'b00011101101000:	sigmoid = 21'b111110011101011110100;
		14'b00011101101001:	sigmoid = 21'b111110011101101010100;
		14'b00011101101010:	sigmoid = 21'b111110011101110110011;
		14'b00011101101011:	sigmoid = 21'b111110011110000010011;
		14'b00011101101100:	sigmoid = 21'b111110011110001110011;
		14'b00011101101101:	sigmoid = 21'b111110011110011010010;
		14'b00011101101110:	sigmoid = 21'b111110011110100110001;
		14'b00011101101111:	sigmoid = 21'b111110011110110010000;
		14'b00011101110000:	sigmoid = 21'b111110011110111101111;
		14'b00011101110001:	sigmoid = 21'b111110011111001001110;
		14'b00011101110010:	sigmoid = 21'b111110011111010101100;
		14'b00011101110011:	sigmoid = 21'b111110011111100001010;
		14'b00011101110100:	sigmoid = 21'b111110011111101101001;
		14'b00011101110101:	sigmoid = 21'b111110011111111000111;
		14'b00011101110110:	sigmoid = 21'b111110100000000100100;
		14'b00011101110111:	sigmoid = 21'b111110100000010000010;
		14'b00011101111000:	sigmoid = 21'b111110100000011011111;
		14'b00011101111001:	sigmoid = 21'b111110100000100111101;
		14'b00011101111010:	sigmoid = 21'b111110100000110011010;
		14'b00011101111011:	sigmoid = 21'b111110100000111110111;
		14'b00011101111100:	sigmoid = 21'b111110100001001010011;
		14'b00011101111101:	sigmoid = 21'b111110100001010110000;
		14'b00011101111110:	sigmoid = 21'b111110100001100001100;
		14'b00011101111111:	sigmoid = 21'b111110100001101101000;
		14'b00011110000000:	sigmoid = 21'b111110100001111000100;
		14'b00011110000001:	sigmoid = 21'b111110100010000100000;
		14'b00011110000010:	sigmoid = 21'b111110100010001111100;
		14'b00011110000011:	sigmoid = 21'b111110100010011011000;
		14'b00011110000100:	sigmoid = 21'b111110100010100110011;
		14'b00011110000101:	sigmoid = 21'b111110100010110001110;
		14'b00011110000110:	sigmoid = 21'b111110100010111101001;
		14'b00011110000111:	sigmoid = 21'b111110100011001000100;
		14'b00011110001000:	sigmoid = 21'b111110100011010011111;
		14'b00011110001001:	sigmoid = 21'b111110100011011111001;
		14'b00011110001010:	sigmoid = 21'b111110100011101010011;
		14'b00011110001011:	sigmoid = 21'b111110100011110101110;
		14'b00011110001100:	sigmoid = 21'b111110100100000001000;
		14'b00011110001101:	sigmoid = 21'b111110100100001100001;
		14'b00011110001110:	sigmoid = 21'b111110100100010111011;
		14'b00011110001111:	sigmoid = 21'b111110100100100010101;
		14'b00011110010000:	sigmoid = 21'b111110100100101101110;
		14'b00011110010001:	sigmoid = 21'b111110100100111000111;
		14'b00011110010010:	sigmoid = 21'b111110100101000100000;
		14'b00011110010011:	sigmoid = 21'b111110100101001111001;
		14'b00011110010100:	sigmoid = 21'b111110100101011010010;
		14'b00011110010101:	sigmoid = 21'b111110100101100101010;
		14'b00011110010110:	sigmoid = 21'b111110100101110000010;
		14'b00011110010111:	sigmoid = 21'b111110100101111011011;
		14'b00011110011000:	sigmoid = 21'b111110100110000110011;
		14'b00011110011001:	sigmoid = 21'b111110100110010001011;
		14'b00011110011010:	sigmoid = 21'b111110100110011100010;
		14'b00011110011011:	sigmoid = 21'b111110100110100111010;
		14'b00011110011100:	sigmoid = 21'b111110100110110010001;
		14'b00011110011101:	sigmoid = 21'b111110100110111101000;
		14'b00011110011110:	sigmoid = 21'b111110100111000111111;
		14'b00011110011111:	sigmoid = 21'b111110100111010010110;
		14'b00011110100000:	sigmoid = 21'b111110100111011101101;
		14'b00011110100001:	sigmoid = 21'b111110100111101000011;
		14'b00011110100010:	sigmoid = 21'b111110100111110011010;
		14'b00011110100011:	sigmoid = 21'b111110100111111110000;
		14'b00011110100100:	sigmoid = 21'b111110101000001000110;
		14'b00011110100101:	sigmoid = 21'b111110101000010011100;
		14'b00011110100110:	sigmoid = 21'b111110101000011110010;
		14'b00011110100111:	sigmoid = 21'b111110101000101000111;
		14'b00011110101000:	sigmoid = 21'b111110101000110011101;
		14'b00011110101001:	sigmoid = 21'b111110101000111110010;
		14'b00011110101010:	sigmoid = 21'b111110101001001000111;
		14'b00011110101011:	sigmoid = 21'b111110101001010011100;
		14'b00011110101100:	sigmoid = 21'b111110101001011110001;
		14'b00011110101101:	sigmoid = 21'b111110101001101000101;
		14'b00011110101110:	sigmoid = 21'b111110101001110011010;
		14'b00011110101111:	sigmoid = 21'b111110101001111101110;
		14'b00011110110000:	sigmoid = 21'b111110101010001000010;
		14'b00011110110001:	sigmoid = 21'b111110101010010010110;
		14'b00011110110010:	sigmoid = 21'b111110101010011101010;
		14'b00011110110011:	sigmoid = 21'b111110101010100111110;
		14'b00011110110100:	sigmoid = 21'b111110101010110010001;
		14'b00011110110101:	sigmoid = 21'b111110101010111100101;
		14'b00011110110110:	sigmoid = 21'b111110101011000111000;
		14'b00011110110111:	sigmoid = 21'b111110101011010001011;
		14'b00011110111000:	sigmoid = 21'b111110101011011011110;
		14'b00011110111001:	sigmoid = 21'b111110101011100110001;
		14'b00011110111010:	sigmoid = 21'b111110101011110000011;
		14'b00011110111011:	sigmoid = 21'b111110101011111010110;
		14'b00011110111100:	sigmoid = 21'b111110101100000101000;
		14'b00011110111101:	sigmoid = 21'b111110101100001111010;
		14'b00011110111110:	sigmoid = 21'b111110101100011001100;
		14'b00011110111111:	sigmoid = 21'b111110101100100011110;
		14'b00011111000000:	sigmoid = 21'b111110101100101101111;
		14'b00011111000001:	sigmoid = 21'b111110101100111000001;
		14'b00011111000010:	sigmoid = 21'b111110101101000010010;
		14'b00011111000011:	sigmoid = 21'b111110101101001100100;
		14'b00011111000100:	sigmoid = 21'b111110101101010110101;
		14'b00011111000101:	sigmoid = 21'b111110101101100000101;
		14'b00011111000110:	sigmoid = 21'b111110101101101010110;
		14'b00011111000111:	sigmoid = 21'b111110101101110100111;
		14'b00011111001000:	sigmoid = 21'b111110101101111110111;
		14'b00011111001001:	sigmoid = 21'b111110101110001001000;
		14'b00011111001010:	sigmoid = 21'b111110101110010011000;
		14'b00011111001011:	sigmoid = 21'b111110101110011101000;
		14'b00011111001100:	sigmoid = 21'b111110101110100111000;
		14'b00011111001101:	sigmoid = 21'b111110101110110000111;
		14'b00011111001110:	sigmoid = 21'b111110101110111010111;
		14'b00011111001111:	sigmoid = 21'b111110101111000100110;
		14'b00011111010000:	sigmoid = 21'b111110101111001110101;
		14'b00011111010001:	sigmoid = 21'b111110101111011000101;
		14'b00011111010010:	sigmoid = 21'b111110101111100010100;
		14'b00011111010011:	sigmoid = 21'b111110101111101100010;
		14'b00011111010100:	sigmoid = 21'b111110101111110110001;
		14'b00011111010101:	sigmoid = 21'b111110110000000000000;
		14'b00011111010110:	sigmoid = 21'b111110110000001001110;
		14'b00011111010111:	sigmoid = 21'b111110110000010011100;
		14'b00011111011000:	sigmoid = 21'b111110110000011101010;
		14'b00011111011001:	sigmoid = 21'b111110110000100111000;
		14'b00011111011010:	sigmoid = 21'b111110110000110000110;
		14'b00011111011011:	sigmoid = 21'b111110110000111010100;
		14'b00011111011100:	sigmoid = 21'b111110110001000100001;
		14'b00011111011101:	sigmoid = 21'b111110110001001101110;
		14'b00011111011110:	sigmoid = 21'b111110110001010111100;
		14'b00011111011111:	sigmoid = 21'b111110110001100001001;
		14'b00011111100000:	sigmoid = 21'b111110110001101010101;
		14'b00011111100001:	sigmoid = 21'b111110110001110100010;
		14'b00011111100010:	sigmoid = 21'b111110110001111101111;
		14'b00011111100011:	sigmoid = 21'b111110110010000111011;
		14'b00011111100100:	sigmoid = 21'b111110110010010001000;
		14'b00011111100101:	sigmoid = 21'b111110110010011010100;
		14'b00011111100110:	sigmoid = 21'b111110110010100100000;
		14'b00011111100111:	sigmoid = 21'b111110110010101101100;
		14'b00011111101000:	sigmoid = 21'b111110110010110111000;
		14'b00011111101001:	sigmoid = 21'b111110110011000000011;
		14'b00011111101010:	sigmoid = 21'b111110110011001001111;
		14'b00011111101011:	sigmoid = 21'b111110110011010011010;
		14'b00011111101100:	sigmoid = 21'b111110110011011100101;
		14'b00011111101101:	sigmoid = 21'b111110110011100110000;
		14'b00011111101110:	sigmoid = 21'b111110110011101111011;
		14'b00011111101111:	sigmoid = 21'b111110110011111000110;
		14'b00011111110000:	sigmoid = 21'b111110110100000010001;
		14'b00011111110001:	sigmoid = 21'b111110110100001011011;
		14'b00011111110010:	sigmoid = 21'b111110110100010100101;
		14'b00011111110011:	sigmoid = 21'b111110110100011110000;
		14'b00011111110100:	sigmoid = 21'b111110110100100111010;
		14'b00011111110101:	sigmoid = 21'b111110110100110000100;
		14'b00011111110110:	sigmoid = 21'b111110110100111001101;
		14'b00011111110111:	sigmoid = 21'b111110110101000010111;
		14'b00011111111000:	sigmoid = 21'b111110110101001100001;
		14'b00011111111001:	sigmoid = 21'b111110110101010101010;
		14'b00011111111010:	sigmoid = 21'b111110110101011110011;
		14'b00011111111011:	sigmoid = 21'b111110110101100111100;
		14'b00011111111100:	sigmoid = 21'b111110110101110000101;
		14'b00011111111101:	sigmoid = 21'b111110110101111001110;
		14'b00011111111110:	sigmoid = 21'b111110110110000010111;
		14'b00011111111111:	sigmoid = 21'b111110110110001011111;
		14'b00100000000000:	sigmoid = 21'b111110110110010101000;
		14'b00100000000001:	sigmoid = 21'b111110110110011110000;
		14'b00100000000010:	sigmoid = 21'b111110110110100111000;
		14'b00100000000011:	sigmoid = 21'b111110110110110000000;
		14'b00100000000100:	sigmoid = 21'b111110110110111001000;
		14'b00100000000101:	sigmoid = 21'b111110110111000010000;
		14'b00100000000110:	sigmoid = 21'b111110110111001010111;
		14'b00100000000111:	sigmoid = 21'b111110110111010011111;
		14'b00100000001000:	sigmoid = 21'b111110110111011100110;
		14'b00100000001001:	sigmoid = 21'b111110110111100101101;
		14'b00100000001010:	sigmoid = 21'b111110110111101110100;
		14'b00100000001011:	sigmoid = 21'b111110110111110111011;
		14'b00100000001100:	sigmoid = 21'b111110111000000000010;
		14'b00100000001101:	sigmoid = 21'b111110111000001001001;
		14'b00100000001110:	sigmoid = 21'b111110111000010001111;
		14'b00100000001111:	sigmoid = 21'b111110111000011010110;
		14'b00100000010000:	sigmoid = 21'b111110111000100011100;
		14'b00100000010001:	sigmoid = 21'b111110111000101100010;
		14'b00100000010010:	sigmoid = 21'b111110111000110101000;
		14'b00100000010011:	sigmoid = 21'b111110111000111101110;
		14'b00100000010100:	sigmoid = 21'b111110111001000110100;
		14'b00100000010101:	sigmoid = 21'b111110111001001111001;
		14'b00100000010110:	sigmoid = 21'b111110111001010111111;
		14'b00100000010111:	sigmoid = 21'b111110111001100000100;
		14'b00100000011000:	sigmoid = 21'b111110111001101001001;
		14'b00100000011001:	sigmoid = 21'b111110111001110001110;
		14'b00100000011010:	sigmoid = 21'b111110111001111010011;
		14'b00100000011011:	sigmoid = 21'b111110111010000011000;
		14'b00100000011100:	sigmoid = 21'b111110111010001011101;
		14'b00100000011101:	sigmoid = 21'b111110111010010100001;
		14'b00100000011110:	sigmoid = 21'b111110111010011100110;
		14'b00100000011111:	sigmoid = 21'b111110111010100101010;
		14'b00100000100000:	sigmoid = 21'b111110111010101101110;
		14'b00100000100001:	sigmoid = 21'b111110111010110110010;
		14'b00100000100010:	sigmoid = 21'b111110111010111110110;
		14'b00100000100011:	sigmoid = 21'b111110111011000111010;
		14'b00100000100100:	sigmoid = 21'b111110111011001111110;
		14'b00100000100101:	sigmoid = 21'b111110111011011000001;
		14'b00100000100110:	sigmoid = 21'b111110111011100000101;
		14'b00100000100111:	sigmoid = 21'b111110111011101001000;
		14'b00100000101000:	sigmoid = 21'b111110111011110001011;
		14'b00100000101001:	sigmoid = 21'b111110111011111001110;
		14'b00100000101010:	sigmoid = 21'b111110111100000010001;
		14'b00100000101011:	sigmoid = 21'b111110111100001010100;
		14'b00100000101100:	sigmoid = 21'b111110111100010010111;
		14'b00100000101101:	sigmoid = 21'b111110111100011011001;
		14'b00100000101110:	sigmoid = 21'b111110111100100011011;
		14'b00100000101111:	sigmoid = 21'b111110111100101011110;
		14'b00100000110000:	sigmoid = 21'b111110111100110100000;
		14'b00100000110001:	sigmoid = 21'b111110111100111100010;
		14'b00100000110010:	sigmoid = 21'b111110111101000100100;
		14'b00100000110011:	sigmoid = 21'b111110111101001100110;
		14'b00100000110100:	sigmoid = 21'b111110111101010100111;
		14'b00100000110101:	sigmoid = 21'b111110111101011101001;
		14'b00100000110110:	sigmoid = 21'b111110111101100101010;
		14'b00100000110111:	sigmoid = 21'b111110111101101101011;
		14'b00100000111000:	sigmoid = 21'b111110111101110101101;
		14'b00100000111001:	sigmoid = 21'b111110111101111101110;
		14'b00100000111010:	sigmoid = 21'b111110111110000101110;
		14'b00100000111011:	sigmoid = 21'b111110111110001101111;
		14'b00100000111100:	sigmoid = 21'b111110111110010110000;
		14'b00100000111101:	sigmoid = 21'b111110111110011110000;
		14'b00100000111110:	sigmoid = 21'b111110111110100110001;
		14'b00100000111111:	sigmoid = 21'b111110111110101110001;
		14'b00100001000000:	sigmoid = 21'b111110111110110110001;
		14'b00100001000001:	sigmoid = 21'b111110111110111110001;
		14'b00100001000010:	sigmoid = 21'b111110111111000110001;
		14'b00100001000011:	sigmoid = 21'b111110111111001110001;
		14'b00100001000100:	sigmoid = 21'b111110111111010110001;
		14'b00100001000101:	sigmoid = 21'b111110111111011110000;
		14'b00100001000110:	sigmoid = 21'b111110111111100110000;
		14'b00100001000111:	sigmoid = 21'b111110111111101101111;
		14'b00100001001000:	sigmoid = 21'b111110111111110101110;
		14'b00100001001001:	sigmoid = 21'b111110111111111101110;
		14'b00100001001010:	sigmoid = 21'b111111000000000101101;
		14'b00100001001011:	sigmoid = 21'b111111000000001101011;
		14'b00100001001100:	sigmoid = 21'b111111000000010101010;
		14'b00100001001101:	sigmoid = 21'b111111000000011101001;
		14'b00100001001110:	sigmoid = 21'b111111000000100100111;
		14'b00100001001111:	sigmoid = 21'b111111000000101100110;
		14'b00100001010000:	sigmoid = 21'b111111000000110100100;
		14'b00100001010001:	sigmoid = 21'b111111000000111100010;
		14'b00100001010010:	sigmoid = 21'b111111000001000100000;
		14'b00100001010011:	sigmoid = 21'b111111000001001011110;
		14'b00100001010100:	sigmoid = 21'b111111000001010011100;
		14'b00100001010101:	sigmoid = 21'b111111000001011011001;
		14'b00100001010110:	sigmoid = 21'b111111000001100010111;
		14'b00100001010111:	sigmoid = 21'b111111000001101010100;
		14'b00100001011000:	sigmoid = 21'b111111000001110010010;
		14'b00100001011001:	sigmoid = 21'b111111000001111001111;
		14'b00100001011010:	sigmoid = 21'b111111000010000001100;
		14'b00100001011011:	sigmoid = 21'b111111000010001001001;
		14'b00100001011100:	sigmoid = 21'b111111000010010000110;
		14'b00100001011101:	sigmoid = 21'b111111000010011000011;
		14'b00100001011110:	sigmoid = 21'b111111000010011111111;
		14'b00100001011111:	sigmoid = 21'b111111000010100111100;
		14'b00100001100000:	sigmoid = 21'b111111000010101111000;
		14'b00100001100001:	sigmoid = 21'b111111000010110110101;
		14'b00100001100010:	sigmoid = 21'b111111000010111110001;
		14'b00100001100011:	sigmoid = 21'b111111000011000101101;
		14'b00100001100100:	sigmoid = 21'b111111000011001101001;
		14'b00100001100101:	sigmoid = 21'b111111000011010100101;
		14'b00100001100110:	sigmoid = 21'b111111000011011100000;
		14'b00100001100111:	sigmoid = 21'b111111000011100011100;
		14'b00100001101000:	sigmoid = 21'b111111000011101010111;
		14'b00100001101001:	sigmoid = 21'b111111000011110010011;
		14'b00100001101010:	sigmoid = 21'b111111000011111001110;
		14'b00100001101011:	sigmoid = 21'b111111000100000001001;
		14'b00100001101100:	sigmoid = 21'b111111000100001000100;
		14'b00100001101101:	sigmoid = 21'b111111000100001111111;
		14'b00100001101110:	sigmoid = 21'b111111000100010111010;
		14'b00100001101111:	sigmoid = 21'b111111000100011110101;
		14'b00100001110000:	sigmoid = 21'b111111000100100101111;
		14'b00100001110001:	sigmoid = 21'b111111000100101101010;
		14'b00100001110010:	sigmoid = 21'b111111000100110100100;
		14'b00100001110011:	sigmoid = 21'b111111000100111011110;
		14'b00100001110100:	sigmoid = 21'b111111000101000011001;
		14'b00100001110101:	sigmoid = 21'b111111000101001010011;
		14'b00100001110110:	sigmoid = 21'b111111000101010001101;
		14'b00100001110111:	sigmoid = 21'b111111000101011000110;
		14'b00100001111000:	sigmoid = 21'b111111000101100000000;
		14'b00100001111001:	sigmoid = 21'b111111000101100111010;
		14'b00100001111010:	sigmoid = 21'b111111000101101110011;
		14'b00100001111011:	sigmoid = 21'b111111000101110101101;
		14'b00100001111100:	sigmoid = 21'b111111000101111100110;
		14'b00100001111101:	sigmoid = 21'b111111000110000011111;
		14'b00100001111110:	sigmoid = 21'b111111000110001011000;
		14'b00100001111111:	sigmoid = 21'b111111000110010010001;
		14'b00100010000000:	sigmoid = 21'b111111000110011001010;
		14'b00100010000001:	sigmoid = 21'b111111000110100000011;
		14'b00100010000010:	sigmoid = 21'b111111000110100111011;
		14'b00100010000011:	sigmoid = 21'b111111000110101110100;
		14'b00100010000100:	sigmoid = 21'b111111000110110101100;
		14'b00100010000101:	sigmoid = 21'b111111000110111100101;
		14'b00100010000110:	sigmoid = 21'b111111000111000011101;
		14'b00100010000111:	sigmoid = 21'b111111000111001010101;
		14'b00100010001000:	sigmoid = 21'b111111000111010001101;
		14'b00100010001001:	sigmoid = 21'b111111000111011000101;
		14'b00100010001010:	sigmoid = 21'b111111000111011111101;
		14'b00100010001011:	sigmoid = 21'b111111000111100110100;
		14'b00100010001100:	sigmoid = 21'b111111000111101101100;
		14'b00100010001101:	sigmoid = 21'b111111000111110100011;
		14'b00100010001110:	sigmoid = 21'b111111000111111011011;
		14'b00100010001111:	sigmoid = 21'b111111001000000010010;
		14'b00100010010000:	sigmoid = 21'b111111001000001001001;
		14'b00100010010001:	sigmoid = 21'b111111001000010000000;
		14'b00100010010010:	sigmoid = 21'b111111001000010110111;
		14'b00100010010011:	sigmoid = 21'b111111001000011101110;
		14'b00100010010100:	sigmoid = 21'b111111001000100100101;
		14'b00100010010101:	sigmoid = 21'b111111001000101011011;
		14'b00100010010110:	sigmoid = 21'b111111001000110010010;
		14'b00100010010111:	sigmoid = 21'b111111001000111001000;
		14'b00100010011000:	sigmoid = 21'b111111001000111111110;
		14'b00100010011001:	sigmoid = 21'b111111001001000110101;
		14'b00100010011010:	sigmoid = 21'b111111001001001101011;
		14'b00100010011011:	sigmoid = 21'b111111001001010100001;
		14'b00100010011100:	sigmoid = 21'b111111001001011010111;
		14'b00100010011101:	sigmoid = 21'b111111001001100001100;
		14'b00100010011110:	sigmoid = 21'b111111001001101000010;
		14'b00100010011111:	sigmoid = 21'b111111001001101111000;
		14'b00100010100000:	sigmoid = 21'b111111001001110101101;
		14'b00100010100001:	sigmoid = 21'b111111001001111100011;
		14'b00100010100010:	sigmoid = 21'b111111001010000011000;
		14'b00100010100011:	sigmoid = 21'b111111001010001001101;
		14'b00100010100100:	sigmoid = 21'b111111001010010000010;
		14'b00100010100101:	sigmoid = 21'b111111001010010110111;
		14'b00100010100110:	sigmoid = 21'b111111001010011101100;
		14'b00100010100111:	sigmoid = 21'b111111001010100100001;
		14'b00100010101000:	sigmoid = 21'b111111001010101010110;
		14'b00100010101001:	sigmoid = 21'b111111001010110001010;
		14'b00100010101010:	sigmoid = 21'b111111001010110111111;
		14'b00100010101011:	sigmoid = 21'b111111001010111110011;
		14'b00100010101100:	sigmoid = 21'b111111001011000100111;
		14'b00100010101101:	sigmoid = 21'b111111001011001011011;
		14'b00100010101110:	sigmoid = 21'b111111001011010010000;
		14'b00100010101111:	sigmoid = 21'b111111001011011000100;
		14'b00100010110000:	sigmoid = 21'b111111001011011110111;
		14'b00100010110001:	sigmoid = 21'b111111001011100101011;
		14'b00100010110010:	sigmoid = 21'b111111001011101011111;
		14'b00100010110011:	sigmoid = 21'b111111001011110010011;
		14'b00100010110100:	sigmoid = 21'b111111001011111000110;
		14'b00100010110101:	sigmoid = 21'b111111001011111111001;
		14'b00100010110110:	sigmoid = 21'b111111001100000101101;
		14'b00100010110111:	sigmoid = 21'b111111001100001100000;
		14'b00100010111000:	sigmoid = 21'b111111001100010010011;
		14'b00100010111001:	sigmoid = 21'b111111001100011000110;
		14'b00100010111010:	sigmoid = 21'b111111001100011111001;
		14'b00100010111011:	sigmoid = 21'b111111001100100101100;
		14'b00100010111100:	sigmoid = 21'b111111001100101011111;
		14'b00100010111101:	sigmoid = 21'b111111001100110010001;
		14'b00100010111110:	sigmoid = 21'b111111001100111000100;
		14'b00100010111111:	sigmoid = 21'b111111001100111110110;
		14'b00100011000000:	sigmoid = 21'b111111001101000101000;
		14'b00100011000001:	sigmoid = 21'b111111001101001011011;
		14'b00100011000010:	sigmoid = 21'b111111001101010001101;
		14'b00100011000011:	sigmoid = 21'b111111001101010111111;
		14'b00100011000100:	sigmoid = 21'b111111001101011110001;
		14'b00100011000101:	sigmoid = 21'b111111001101100100011;
		14'b00100011000110:	sigmoid = 21'b111111001101101010100;
		14'b00100011000111:	sigmoid = 21'b111111001101110000110;
		14'b00100011001000:	sigmoid = 21'b111111001101110111000;
		14'b00100011001001:	sigmoid = 21'b111111001101111101001;
		14'b00100011001010:	sigmoid = 21'b111111001110000011011;
		14'b00100011001011:	sigmoid = 21'b111111001110001001100;
		14'b00100011001100:	sigmoid = 21'b111111001110001111101;
		14'b00100011001101:	sigmoid = 21'b111111001110010101110;
		14'b00100011001110:	sigmoid = 21'b111111001110011011111;
		14'b00100011001111:	sigmoid = 21'b111111001110100010000;
		14'b00100011010000:	sigmoid = 21'b111111001110101000001;
		14'b00100011010001:	sigmoid = 21'b111111001110101110010;
		14'b00100011010010:	sigmoid = 21'b111111001110110100010;
		14'b00100011010011:	sigmoid = 21'b111111001110111010011;
		14'b00100011010100:	sigmoid = 21'b111111001111000000011;
		14'b00100011010101:	sigmoid = 21'b111111001111000110100;
		14'b00100011010110:	sigmoid = 21'b111111001111001100100;
		14'b00100011010111:	sigmoid = 21'b111111001111010010100;
		14'b00100011011000:	sigmoid = 21'b111111001111011000100;
		14'b00100011011001:	sigmoid = 21'b111111001111011110100;
		14'b00100011011010:	sigmoid = 21'b111111001111100100100;
		14'b00100011011011:	sigmoid = 21'b111111001111101010100;
		14'b00100011011100:	sigmoid = 21'b111111001111110000100;
		14'b00100011011101:	sigmoid = 21'b111111001111110110011;
		14'b00100011011110:	sigmoid = 21'b111111001111111100011;
		14'b00100011011111:	sigmoid = 21'b111111010000000010010;
		14'b00100011100000:	sigmoid = 21'b111111010000001000010;
		14'b00100011100001:	sigmoid = 21'b111111010000001110001;
		14'b00100011100010:	sigmoid = 21'b111111010000010100000;
		14'b00100011100011:	sigmoid = 21'b111111010000011001111;
		14'b00100011100100:	sigmoid = 21'b111111010000011111110;
		14'b00100011100101:	sigmoid = 21'b111111010000100101101;
		14'b00100011100110:	sigmoid = 21'b111111010000101011100;
		14'b00100011100111:	sigmoid = 21'b111111010000110001011;
		14'b00100011101000:	sigmoid = 21'b111111010000110111001;
		14'b00100011101001:	sigmoid = 21'b111111010000111101000;
		14'b00100011101010:	sigmoid = 21'b111111010001000010110;
		14'b00100011101011:	sigmoid = 21'b111111010001001000101;
		14'b00100011101100:	sigmoid = 21'b111111010001001110011;
		14'b00100011101101:	sigmoid = 21'b111111010001010100001;
		14'b00100011101110:	sigmoid = 21'b111111010001011001111;
		14'b00100011101111:	sigmoid = 21'b111111010001011111101;
		14'b00100011110000:	sigmoid = 21'b111111010001100101011;
		14'b00100011110001:	sigmoid = 21'b111111010001101011001;
		14'b00100011110010:	sigmoid = 21'b111111010001110000111;
		14'b00100011110011:	sigmoid = 21'b111111010001110110100;
		14'b00100011110100:	sigmoid = 21'b111111010001111100010;
		14'b00100011110101:	sigmoid = 21'b111111010010000001111;
		14'b00100011110110:	sigmoid = 21'b111111010010000111101;
		14'b00100011110111:	sigmoid = 21'b111111010010001101010;
		14'b00100011111000:	sigmoid = 21'b111111010010010010111;
		14'b00100011111001:	sigmoid = 21'b111111010010011000101;
		14'b00100011111010:	sigmoid = 21'b111111010010011110010;
		14'b00100011111011:	sigmoid = 21'b111111010010100011111;
		14'b00100011111100:	sigmoid = 21'b111111010010101001011;
		14'b00100011111101:	sigmoid = 21'b111111010010101111000;
		14'b00100011111110:	sigmoid = 21'b111111010010110100101;
		14'b00100011111111:	sigmoid = 21'b111111010010111010010;
		14'b00100100000000:	sigmoid = 21'b111111010010111111110;
		14'b00100100000001:	sigmoid = 21'b111111010011000101011;
		14'b00100100000010:	sigmoid = 21'b111111010011001010111;
		14'b00100100000011:	sigmoid = 21'b111111010011010000011;
		14'b00100100000100:	sigmoid = 21'b111111010011010110000;
		14'b00100100000101:	sigmoid = 21'b111111010011011011100;
		14'b00100100000110:	sigmoid = 21'b111111010011100001000;
		14'b00100100000111:	sigmoid = 21'b111111010011100110100;
		14'b00100100001000:	sigmoid = 21'b111111010011101100000;
		14'b00100100001001:	sigmoid = 21'b111111010011110001011;
		14'b00100100001010:	sigmoid = 21'b111111010011110110111;
		14'b00100100001011:	sigmoid = 21'b111111010011111100011;
		14'b00100100001100:	sigmoid = 21'b111111010100000001110;
		14'b00100100001101:	sigmoid = 21'b111111010100000111010;
		14'b00100100001110:	sigmoid = 21'b111111010100001100101;
		14'b00100100001111:	sigmoid = 21'b111111010100010010000;
		14'b00100100010000:	sigmoid = 21'b111111010100010111100;
		14'b00100100010001:	sigmoid = 21'b111111010100011100111;
		14'b00100100010010:	sigmoid = 21'b111111010100100010010;
		14'b00100100010011:	sigmoid = 21'b111111010100100111101;
		14'b00100100010100:	sigmoid = 21'b111111010100101101000;
		14'b00100100010101:	sigmoid = 21'b111111010100110010010;
		14'b00100100010110:	sigmoid = 21'b111111010100110111101;
		14'b00100100010111:	sigmoid = 21'b111111010100111101000;
		14'b00100100011000:	sigmoid = 21'b111111010101000010010;
		14'b00100100011001:	sigmoid = 21'b111111010101000111101;
		14'b00100100011010:	sigmoid = 21'b111111010101001100111;
		14'b00100100011011:	sigmoid = 21'b111111010101010010001;
		14'b00100100011100:	sigmoid = 21'b111111010101010111100;
		14'b00100100011101:	sigmoid = 21'b111111010101011100110;
		14'b00100100011110:	sigmoid = 21'b111111010101100010000;
		14'b00100100011111:	sigmoid = 21'b111111010101100111010;
		14'b00100100100000:	sigmoid = 21'b111111010101101100100;
		14'b00100100100001:	sigmoid = 21'b111111010101110001110;
		14'b00100100100010:	sigmoid = 21'b111111010101110110111;
		14'b00100100100011:	sigmoid = 21'b111111010101111100001;
		14'b00100100100100:	sigmoid = 21'b111111010110000001011;
		14'b00100100100101:	sigmoid = 21'b111111010110000110100;
		14'b00100100100110:	sigmoid = 21'b111111010110001011110;
		14'b00100100100111:	sigmoid = 21'b111111010110010000111;
		14'b00100100101000:	sigmoid = 21'b111111010110010110000;
		14'b00100100101001:	sigmoid = 21'b111111010110011011001;
		14'b00100100101010:	sigmoid = 21'b111111010110100000010;
		14'b00100100101011:	sigmoid = 21'b111111010110100101100;
		14'b00100100101100:	sigmoid = 21'b111111010110101010100;
		14'b00100100101101:	sigmoid = 21'b111111010110101111101;
		14'b00100100101110:	sigmoid = 21'b111111010110110100110;
		14'b00100100101111:	sigmoid = 21'b111111010110111001111;
		14'b00100100110000:	sigmoid = 21'b111111010110111111000;
		14'b00100100110001:	sigmoid = 21'b111111010111000100000;
		14'b00100100110010:	sigmoid = 21'b111111010111001001001;
		14'b00100100110011:	sigmoid = 21'b111111010111001110001;
		14'b00100100110100:	sigmoid = 21'b111111010111010011001;
		14'b00100100110101:	sigmoid = 21'b111111010111011000010;
		14'b00100100110110:	sigmoid = 21'b111111010111011101010;
		14'b00100100110111:	sigmoid = 21'b111111010111100010010;
		14'b00100100111000:	sigmoid = 21'b111111010111100111010;
		14'b00100100111001:	sigmoid = 21'b111111010111101100010;
		14'b00100100111010:	sigmoid = 21'b111111010111110001010;
		14'b00100100111011:	sigmoid = 21'b111111010111110110010;
		14'b00100100111100:	sigmoid = 21'b111111010111111011001;
		14'b00100100111101:	sigmoid = 21'b111111011000000000001;
		14'b00100100111110:	sigmoid = 21'b111111011000000101000;
		14'b00100100111111:	sigmoid = 21'b111111011000001010000;
		14'b00100101000000:	sigmoid = 21'b111111011000001110111;
		14'b00100101000001:	sigmoid = 21'b111111011000010011111;
		14'b00100101000010:	sigmoid = 21'b111111011000011000110;
		14'b00100101000011:	sigmoid = 21'b111111011000011101101;
		14'b00100101000100:	sigmoid = 21'b111111011000100010100;
		14'b00100101000101:	sigmoid = 21'b111111011000100111011;
		14'b00100101000110:	sigmoid = 21'b111111011000101100010;
		14'b00100101000111:	sigmoid = 21'b111111011000110001001;
		14'b00100101001000:	sigmoid = 21'b111111011000110110000;
		14'b00100101001001:	sigmoid = 21'b111111011000111010111;
		14'b00100101001010:	sigmoid = 21'b111111011000111111101;
		14'b00100101001011:	sigmoid = 21'b111111011001000100100;
		14'b00100101001100:	sigmoid = 21'b111111011001001001011;
		14'b00100101001101:	sigmoid = 21'b111111011001001110001;
		14'b00100101001110:	sigmoid = 21'b111111011001010010111;
		14'b00100101001111:	sigmoid = 21'b111111011001010111110;
		14'b00100101010000:	sigmoid = 21'b111111011001011100100;
		14'b00100101010001:	sigmoid = 21'b111111011001100001010;
		14'b00100101010010:	sigmoid = 21'b111111011001100110000;
		14'b00100101010011:	sigmoid = 21'b111111011001101010110;
		14'b00100101010100:	sigmoid = 21'b111111011001101111100;
		14'b00100101010101:	sigmoid = 21'b111111011001110100010;
		14'b00100101010110:	sigmoid = 21'b111111011001111001000;
		14'b00100101010111:	sigmoid = 21'b111111011001111101101;
		14'b00100101011000:	sigmoid = 21'b111111011010000010011;
		14'b00100101011001:	sigmoid = 21'b111111011010000111001;
		14'b00100101011010:	sigmoid = 21'b111111011010001011110;
		14'b00100101011011:	sigmoid = 21'b111111011010010000100;
		14'b00100101011100:	sigmoid = 21'b111111011010010101001;
		14'b00100101011101:	sigmoid = 21'b111111011010011001110;
		14'b00100101011110:	sigmoid = 21'b111111011010011110011;
		14'b00100101011111:	sigmoid = 21'b111111011010100011001;
		14'b00100101100000:	sigmoid = 21'b111111011010100111110;
		14'b00100101100001:	sigmoid = 21'b111111011010101100011;
		14'b00100101100010:	sigmoid = 21'b111111011010110001000;
		14'b00100101100011:	sigmoid = 21'b111111011010110101100;
		14'b00100101100100:	sigmoid = 21'b111111011010111010001;
		14'b00100101100101:	sigmoid = 21'b111111011010111110110;
		14'b00100101100110:	sigmoid = 21'b111111011011000011011;
		14'b00100101100111:	sigmoid = 21'b111111011011000111111;
		14'b00100101101000:	sigmoid = 21'b111111011011001100100;
		14'b00100101101001:	sigmoid = 21'b111111011011010001000;
		14'b00100101101010:	sigmoid = 21'b111111011011010101100;
		14'b00100101101011:	sigmoid = 21'b111111011011011010001;
		14'b00100101101100:	sigmoid = 21'b111111011011011110101;
		14'b00100101101101:	sigmoid = 21'b111111011011100011001;
		14'b00100101101110:	sigmoid = 21'b111111011011100111101;
		14'b00100101101111:	sigmoid = 21'b111111011011101100001;
		14'b00100101110000:	sigmoid = 21'b111111011011110000101;
		14'b00100101110001:	sigmoid = 21'b111111011011110101001;
		14'b00100101110010:	sigmoid = 21'b111111011011111001101;
		14'b00100101110011:	sigmoid = 21'b111111011011111110001;
		14'b00100101110100:	sigmoid = 21'b111111011100000010100;
		14'b00100101110101:	sigmoid = 21'b111111011100000111000;
		14'b00100101110110:	sigmoid = 21'b111111011100001011100;
		14'b00100101110111:	sigmoid = 21'b111111011100001111111;
		14'b00100101111000:	sigmoid = 21'b111111011100010100010;
		14'b00100101111001:	sigmoid = 21'b111111011100011000110;
		14'b00100101111010:	sigmoid = 21'b111111011100011101001;
		14'b00100101111011:	sigmoid = 21'b111111011100100001100;
		14'b00100101111100:	sigmoid = 21'b111111011100100101111;
		14'b00100101111101:	sigmoid = 21'b111111011100101010010;
		14'b00100101111110:	sigmoid = 21'b111111011100101110101;
		14'b00100101111111:	sigmoid = 21'b111111011100110011000;
		14'b00100110000000:	sigmoid = 21'b111111011100110111011;
		14'b00100110000001:	sigmoid = 21'b111111011100111011110;
		14'b00100110000010:	sigmoid = 21'b111111011101000000001;
		14'b00100110000011:	sigmoid = 21'b111111011101000100011;
		14'b00100110000100:	sigmoid = 21'b111111011101001000110;
		14'b00100110000101:	sigmoid = 21'b111111011101001101001;
		14'b00100110000110:	sigmoid = 21'b111111011101010001011;
		14'b00100110000111:	sigmoid = 21'b111111011101010101101;
		14'b00100110001000:	sigmoid = 21'b111111011101011010000;
		14'b00100110001001:	sigmoid = 21'b111111011101011110010;
		14'b00100110001010:	sigmoid = 21'b111111011101100010100;
		14'b00100110001011:	sigmoid = 21'b111111011101100110110;
		14'b00100110001100:	sigmoid = 21'b111111011101101011000;
		14'b00100110001101:	sigmoid = 21'b111111011101101111010;
		14'b00100110001110:	sigmoid = 21'b111111011101110011100;
		14'b00100110001111:	sigmoid = 21'b111111011101110111110;
		14'b00100110010000:	sigmoid = 21'b111111011101111100000;
		14'b00100110010001:	sigmoid = 21'b111111011110000000010;
		14'b00100110010010:	sigmoid = 21'b111111011110000100011;
		14'b00100110010011:	sigmoid = 21'b111111011110001000101;
		14'b00100110010100:	sigmoid = 21'b111111011110001100111;
		14'b00100110010101:	sigmoid = 21'b111111011110010001000;
		14'b00100110010110:	sigmoid = 21'b111111011110010101010;
		14'b00100110010111:	sigmoid = 21'b111111011110011001011;
		14'b00100110011000:	sigmoid = 21'b111111011110011101100;
		14'b00100110011001:	sigmoid = 21'b111111011110100001101;
		14'b00100110011010:	sigmoid = 21'b111111011110100101111;
		14'b00100110011011:	sigmoid = 21'b111111011110101010000;
		14'b00100110011100:	sigmoid = 21'b111111011110101110001;
		14'b00100110011101:	sigmoid = 21'b111111011110110010010;
		14'b00100110011110:	sigmoid = 21'b111111011110110110011;
		14'b00100110011111:	sigmoid = 21'b111111011110111010011;
		14'b00100110100000:	sigmoid = 21'b111111011110111110100;
		14'b00100110100001:	sigmoid = 21'b111111011111000010101;
		14'b00100110100010:	sigmoid = 21'b111111011111000110110;
		14'b00100110100011:	sigmoid = 21'b111111011111001010110;
		14'b00100110100100:	sigmoid = 21'b111111011111001110111;
		14'b00100110100101:	sigmoid = 21'b111111011111010010111;
		14'b00100110100110:	sigmoid = 21'b111111011111010111000;
		14'b00100110100111:	sigmoid = 21'b111111011111011011000;
		14'b00100110101000:	sigmoid = 21'b111111011111011111000;
		14'b00100110101001:	sigmoid = 21'b111111011111100011001;
		14'b00100110101010:	sigmoid = 21'b111111011111100111001;
		14'b00100110101011:	sigmoid = 21'b111111011111101011001;
		14'b00100110101100:	sigmoid = 21'b111111011111101111001;
		14'b00100110101101:	sigmoid = 21'b111111011111110011001;
		14'b00100110101110:	sigmoid = 21'b111111011111110111001;
		14'b00100110101111:	sigmoid = 21'b111111011111111011001;
		14'b00100110110000:	sigmoid = 21'b111111011111111111000;
		14'b00100110110001:	sigmoid = 21'b111111100000000011000;
		14'b00100110110010:	sigmoid = 21'b111111100000000111000;
		14'b00100110110011:	sigmoid = 21'b111111100000001010111;
		14'b00100110110100:	sigmoid = 21'b111111100000001110111;
		14'b00100110110101:	sigmoid = 21'b111111100000010010110;
		14'b00100110110110:	sigmoid = 21'b111111100000010110110;
		14'b00100110110111:	sigmoid = 21'b111111100000011010101;
		14'b00100110111000:	sigmoid = 21'b111111100000011110101;
		14'b00100110111001:	sigmoid = 21'b111111100000100010100;
		14'b00100110111010:	sigmoid = 21'b111111100000100110011;
		14'b00100110111011:	sigmoid = 21'b111111100000101010010;
		14'b00100110111100:	sigmoid = 21'b111111100000101110001;
		14'b00100110111101:	sigmoid = 21'b111111100000110010000;
		14'b00100110111110:	sigmoid = 21'b111111100000110101111;
		14'b00100110111111:	sigmoid = 21'b111111100000111001110;
		14'b00100111000000:	sigmoid = 21'b111111100000111101101;
		14'b00100111000001:	sigmoid = 21'b111111100001000001100;
		14'b00100111000010:	sigmoid = 21'b111111100001000101010;
		14'b00100111000011:	sigmoid = 21'b111111100001001001001;
		14'b00100111000100:	sigmoid = 21'b111111100001001101000;
		14'b00100111000101:	sigmoid = 21'b111111100001010000110;
		14'b00100111000110:	sigmoid = 21'b111111100001010100101;
		14'b00100111000111:	sigmoid = 21'b111111100001011000011;
		14'b00100111001000:	sigmoid = 21'b111111100001011100001;
		14'b00100111001001:	sigmoid = 21'b111111100001100000000;
		14'b00100111001010:	sigmoid = 21'b111111100001100011110;
		14'b00100111001011:	sigmoid = 21'b111111100001100111100;
		14'b00100111001100:	sigmoid = 21'b111111100001101011010;
		14'b00100111001101:	sigmoid = 21'b111111100001101111000;
		14'b00100111001110:	sigmoid = 21'b111111100001110010110;
		14'b00100111001111:	sigmoid = 21'b111111100001110110100;
		14'b00100111010000:	sigmoid = 21'b111111100001111010010;
		14'b00100111010001:	sigmoid = 21'b111111100001111110000;
		14'b00100111010010:	sigmoid = 21'b111111100010000001110;
		14'b00100111010011:	sigmoid = 21'b111111100010000101100;
		14'b00100111010100:	sigmoid = 21'b111111100010001001001;
		14'b00100111010101:	sigmoid = 21'b111111100010001100111;
		14'b00100111010110:	sigmoid = 21'b111111100010010000100;
		14'b00100111010111:	sigmoid = 21'b111111100010010100010;
		14'b00100111011000:	sigmoid = 21'b111111100010010111111;
		14'b00100111011001:	sigmoid = 21'b111111100010011011101;
		14'b00100111011010:	sigmoid = 21'b111111100010011111010;
		14'b00100111011011:	sigmoid = 21'b111111100010100010111;
		14'b00100111011100:	sigmoid = 21'b111111100010100110100;
		14'b00100111011101:	sigmoid = 21'b111111100010101010010;
		14'b00100111011110:	sigmoid = 21'b111111100010101101111;
		14'b00100111011111:	sigmoid = 21'b111111100010110001100;
		14'b00100111100000:	sigmoid = 21'b111111100010110101001;
		14'b00100111100001:	sigmoid = 21'b111111100010111000110;
		14'b00100111100010:	sigmoid = 21'b111111100010111100011;
		14'b00100111100011:	sigmoid = 21'b111111100010111111111;
		14'b00100111100100:	sigmoid = 21'b111111100011000011100;
		14'b00100111100101:	sigmoid = 21'b111111100011000111001;
		14'b00100111100110:	sigmoid = 21'b111111100011001010110;
		14'b00100111100111:	sigmoid = 21'b111111100011001110010;
		14'b00100111101000:	sigmoid = 21'b111111100011010001111;
		14'b00100111101001:	sigmoid = 21'b111111100011010101011;
		14'b00100111101010:	sigmoid = 21'b111111100011011001000;
		14'b00100111101011:	sigmoid = 21'b111111100011011100100;
		14'b00100111101100:	sigmoid = 21'b111111100011100000000;
		14'b00100111101101:	sigmoid = 21'b111111100011100011101;
		14'b00100111101110:	sigmoid = 21'b111111100011100111001;
		14'b00100111101111:	sigmoid = 21'b111111100011101010101;
		14'b00100111110000:	sigmoid = 21'b111111100011101110001;
		14'b00100111110001:	sigmoid = 21'b111111100011110001101;
		14'b00100111110010:	sigmoid = 21'b111111100011110101001;
		14'b00100111110011:	sigmoid = 21'b111111100011111000101;
		14'b00100111110100:	sigmoid = 21'b111111100011111100001;
		14'b00100111110101:	sigmoid = 21'b111111100011111111101;
		14'b00100111110110:	sigmoid = 21'b111111100100000011001;
		14'b00100111110111:	sigmoid = 21'b111111100100000110100;
		14'b00100111111000:	sigmoid = 21'b111111100100001010000;
		14'b00100111111001:	sigmoid = 21'b111111100100001101100;
		14'b00100111111010:	sigmoid = 21'b111111100100010000111;
		14'b00100111111011:	sigmoid = 21'b111111100100010100011;
		14'b00100111111100:	sigmoid = 21'b111111100100010111110;
		14'b00100111111101:	sigmoid = 21'b111111100100011011010;
		14'b00100111111110:	sigmoid = 21'b111111100100011110101;
		14'b00100111111111:	sigmoid = 21'b111111100100100010000;
		14'b00101000000000:	sigmoid = 21'b111111100100100101100;
		14'b00101000000001:	sigmoid = 21'b111111100100101000111;
		14'b00101000000010:	sigmoid = 21'b111111100100101100010;
		14'b00101000000011:	sigmoid = 21'b111111100100101111101;
		14'b00101000000100:	sigmoid = 21'b111111100100110011000;
		14'b00101000000101:	sigmoid = 21'b111111100100110110011;
		14'b00101000000110:	sigmoid = 21'b111111100100111001110;
		14'b00101000000111:	sigmoid = 21'b111111100100111101001;
		14'b00101000001000:	sigmoid = 21'b111111100101000000100;
		14'b00101000001001:	sigmoid = 21'b111111100101000011111;
		14'b00101000001010:	sigmoid = 21'b111111100101000111001;
		14'b00101000001011:	sigmoid = 21'b111111100101001010100;
		14'b00101000001100:	sigmoid = 21'b111111100101001101111;
		14'b00101000001101:	sigmoid = 21'b111111100101010001001;
		14'b00101000001110:	sigmoid = 21'b111111100101010100100;
		14'b00101000001111:	sigmoid = 21'b111111100101010111110;
		14'b00101000010000:	sigmoid = 21'b111111100101011011001;
		14'b00101000010001:	sigmoid = 21'b111111100101011110011;
		14'b00101000010010:	sigmoid = 21'b111111100101100001101;
		14'b00101000010011:	sigmoid = 21'b111111100101100101000;
		14'b00101000010100:	sigmoid = 21'b111111100101101000010;
		14'b00101000010101:	sigmoid = 21'b111111100101101011100;
		14'b00101000010110:	sigmoid = 21'b111111100101101110110;
		14'b00101000010111:	sigmoid = 21'b111111100101110010000;
		14'b00101000011000:	sigmoid = 21'b111111100101110101010;
		14'b00101000011001:	sigmoid = 21'b111111100101111000100;
		14'b00101000011010:	sigmoid = 21'b111111100101111011110;
		14'b00101000011011:	sigmoid = 21'b111111100101111111000;
		14'b00101000011100:	sigmoid = 21'b111111100110000010010;
		14'b00101000011101:	sigmoid = 21'b111111100110000101100;
		14'b00101000011110:	sigmoid = 21'b111111100110001000101;
		14'b00101000011111:	sigmoid = 21'b111111100110001011111;
		14'b00101000100000:	sigmoid = 21'b111111100110001111001;
		14'b00101000100001:	sigmoid = 21'b111111100110010010010;
		14'b00101000100010:	sigmoid = 21'b111111100110010101100;
		14'b00101000100011:	sigmoid = 21'b111111100110011000101;
		14'b00101000100100:	sigmoid = 21'b111111100110011011111;
		14'b00101000100101:	sigmoid = 21'b111111100110011111000;
		14'b00101000100110:	sigmoid = 21'b111111100110100010001;
		14'b00101000100111:	sigmoid = 21'b111111100110100101011;
		14'b00101000101000:	sigmoid = 21'b111111100110101000100;
		14'b00101000101001:	sigmoid = 21'b111111100110101011101;
		14'b00101000101010:	sigmoid = 21'b111111100110101110110;
		14'b00101000101011:	sigmoid = 21'b111111100110110001111;
		14'b00101000101100:	sigmoid = 21'b111111100110110101000;
		14'b00101000101101:	sigmoid = 21'b111111100110111000001;
		14'b00101000101110:	sigmoid = 21'b111111100110111011010;
		14'b00101000101111:	sigmoid = 21'b111111100110111110011;
		14'b00101000110000:	sigmoid = 21'b111111100111000001100;
		14'b00101000110001:	sigmoid = 21'b111111100111000100101;
		14'b00101000110010:	sigmoid = 21'b111111100111000111110;
		14'b00101000110011:	sigmoid = 21'b111111100111001010110;
		14'b00101000110100:	sigmoid = 21'b111111100111001101111;
		14'b00101000110101:	sigmoid = 21'b111111100111010001000;
		14'b00101000110110:	sigmoid = 21'b111111100111010100000;
		14'b00101000110111:	sigmoid = 21'b111111100111010111001;
		14'b00101000111000:	sigmoid = 21'b111111100111011010001;
		14'b00101000111001:	sigmoid = 21'b111111100111011101001;
		14'b00101000111010:	sigmoid = 21'b111111100111100000010;
		14'b00101000111011:	sigmoid = 21'b111111100111100011010;
		14'b00101000111100:	sigmoid = 21'b111111100111100110010;
		14'b00101000111101:	sigmoid = 21'b111111100111101001011;
		14'b00101000111110:	sigmoid = 21'b111111100111101100011;
		14'b00101000111111:	sigmoid = 21'b111111100111101111011;
		14'b00101001000000:	sigmoid = 21'b111111100111110010011;
		14'b00101001000001:	sigmoid = 21'b111111100111110101011;
		14'b00101001000010:	sigmoid = 21'b111111100111111000011;
		14'b00101001000011:	sigmoid = 21'b111111100111111011011;
		14'b00101001000100:	sigmoid = 21'b111111100111111110011;
		14'b00101001000101:	sigmoid = 21'b111111101000000001011;
		14'b00101001000110:	sigmoid = 21'b111111101000000100011;
		14'b00101001000111:	sigmoid = 21'b111111101000000111010;
		14'b00101001001000:	sigmoid = 21'b111111101000001010010;
		14'b00101001001001:	sigmoid = 21'b111111101000001101010;
		14'b00101001001010:	sigmoid = 21'b111111101000010000001;
		14'b00101001001011:	sigmoid = 21'b111111101000010011001;
		14'b00101001001100:	sigmoid = 21'b111111101000010110001;
		14'b00101001001101:	sigmoid = 21'b111111101000011001000;
		14'b00101001001110:	sigmoid = 21'b111111101000011100000;
		14'b00101001001111:	sigmoid = 21'b111111101000011110111;
		14'b00101001010000:	sigmoid = 21'b111111101000100001110;
		14'b00101001010001:	sigmoid = 21'b111111101000100100110;
		14'b00101001010010:	sigmoid = 21'b111111101000100111101;
		14'b00101001010011:	sigmoid = 21'b111111101000101010100;
		14'b00101001010100:	sigmoid = 21'b111111101000101101011;
		14'b00101001010101:	sigmoid = 21'b111111101000110000010;
		14'b00101001010110:	sigmoid = 21'b111111101000110011010;
		14'b00101001010111:	sigmoid = 21'b111111101000110110001;
		14'b00101001011000:	sigmoid = 21'b111111101000111001000;
		14'b00101001011001:	sigmoid = 21'b111111101000111011111;
		14'b00101001011010:	sigmoid = 21'b111111101000111110101;
		14'b00101001011011:	sigmoid = 21'b111111101001000001100;
		14'b00101001011100:	sigmoid = 21'b111111101001000100011;
		14'b00101001011101:	sigmoid = 21'b111111101001000111010;
		14'b00101001011110:	sigmoid = 21'b111111101001001010001;
		14'b00101001011111:	sigmoid = 21'b111111101001001100111;
		14'b00101001100000:	sigmoid = 21'b111111101001001111110;
		14'b00101001100001:	sigmoid = 21'b111111101001010010101;
		14'b00101001100010:	sigmoid = 21'b111111101001010101011;
		14'b00101001100011:	sigmoid = 21'b111111101001011000010;
		14'b00101001100100:	sigmoid = 21'b111111101001011011000;
		14'b00101001100101:	sigmoid = 21'b111111101001011101111;
		14'b00101001100110:	sigmoid = 21'b111111101001100000101;
		14'b00101001100111:	sigmoid = 21'b111111101001100011011;
		14'b00101001101000:	sigmoid = 21'b111111101001100110010;
		14'b00101001101001:	sigmoid = 21'b111111101001101001000;
		14'b00101001101010:	sigmoid = 21'b111111101001101011110;
		14'b00101001101011:	sigmoid = 21'b111111101001101110100;
		14'b00101001101100:	sigmoid = 21'b111111101001110001010;
		14'b00101001101101:	sigmoid = 21'b111111101001110100000;
		14'b00101001101110:	sigmoid = 21'b111111101001110110111;
		14'b00101001101111:	sigmoid = 21'b111111101001111001101;
		14'b00101001110000:	sigmoid = 21'b111111101001111100010;
		14'b00101001110001:	sigmoid = 21'b111111101001111111000;
		14'b00101001110010:	sigmoid = 21'b111111101010000001110;
		14'b00101001110011:	sigmoid = 21'b111111101010000100100;
		14'b00101001110100:	sigmoid = 21'b111111101010000111010;
		14'b00101001110101:	sigmoid = 21'b111111101010001010000;
		14'b00101001110110:	sigmoid = 21'b111111101010001100101;
		14'b00101001110111:	sigmoid = 21'b111111101010001111011;
		14'b00101001111000:	sigmoid = 21'b111111101010010010001;
		14'b00101001111001:	sigmoid = 21'b111111101010010100110;
		14'b00101001111010:	sigmoid = 21'b111111101010010111100;
		14'b00101001111011:	sigmoid = 21'b111111101010011010001;
		14'b00101001111100:	sigmoid = 21'b111111101010011100111;
		14'b00101001111101:	sigmoid = 21'b111111101010011111100;
		14'b00101001111110:	sigmoid = 21'b111111101010100010001;
		14'b00101001111111:	sigmoid = 21'b111111101010100100111;
		14'b00101010000000:	sigmoid = 21'b111111101010100111100;
		14'b00101010000001:	sigmoid = 21'b111111101010101010001;
		14'b00101010000010:	sigmoid = 21'b111111101010101100111;
		14'b00101010000011:	sigmoid = 21'b111111101010101111100;
		14'b00101010000100:	sigmoid = 21'b111111101010110010001;
		14'b00101010000101:	sigmoid = 21'b111111101010110100110;
		14'b00101010000110:	sigmoid = 21'b111111101010110111011;
		14'b00101010000111:	sigmoid = 21'b111111101010111010000;
		14'b00101010001000:	sigmoid = 21'b111111101010111100101;
		14'b00101010001001:	sigmoid = 21'b111111101010111111010;
		14'b00101010001010:	sigmoid = 21'b111111101011000001111;
		14'b00101010001011:	sigmoid = 21'b111111101011000100100;
		14'b00101010001100:	sigmoid = 21'b111111101011000111000;
		14'b00101010001101:	sigmoid = 21'b111111101011001001101;
		14'b00101010001110:	sigmoid = 21'b111111101011001100010;
		14'b00101010001111:	sigmoid = 21'b111111101011001110111;
		14'b00101010010000:	sigmoid = 21'b111111101011010001011;
		14'b00101010010001:	sigmoid = 21'b111111101011010100000;
		14'b00101010010010:	sigmoid = 21'b111111101011010110100;
		14'b00101010010011:	sigmoid = 21'b111111101011011001001;
		14'b00101010010100:	sigmoid = 21'b111111101011011011101;
		14'b00101010010101:	sigmoid = 21'b111111101011011110010;
		14'b00101010010110:	sigmoid = 21'b111111101011100000110;
		14'b00101010010111:	sigmoid = 21'b111111101011100011011;
		14'b00101010011000:	sigmoid = 21'b111111101011100101111;
		14'b00101010011001:	sigmoid = 21'b111111101011101000011;
		14'b00101010011010:	sigmoid = 21'b111111101011101010111;
		14'b00101010011011:	sigmoid = 21'b111111101011101101100;
		14'b00101010011100:	sigmoid = 21'b111111101011110000000;
		14'b00101010011101:	sigmoid = 21'b111111101011110010100;
		14'b00101010011110:	sigmoid = 21'b111111101011110101000;
		14'b00101010011111:	sigmoid = 21'b111111101011110111100;
		14'b00101010100000:	sigmoid = 21'b111111101011111010000;
		14'b00101010100001:	sigmoid = 21'b111111101011111100100;
		14'b00101010100010:	sigmoid = 21'b111111101011111111000;
		14'b00101010100011:	sigmoid = 21'b111111101100000001100;
		14'b00101010100100:	sigmoid = 21'b111111101100000100000;
		14'b00101010100101:	sigmoid = 21'b111111101100000110100;
		14'b00101010100110:	sigmoid = 21'b111111101100001000111;
		14'b00101010100111:	sigmoid = 21'b111111101100001011011;
		14'b00101010101000:	sigmoid = 21'b111111101100001101111;
		14'b00101010101001:	sigmoid = 21'b111111101100010000011;
		14'b00101010101010:	sigmoid = 21'b111111101100010010110;
		14'b00101010101011:	sigmoid = 21'b111111101100010101010;
		14'b00101010101100:	sigmoid = 21'b111111101100010111101;
		14'b00101010101101:	sigmoid = 21'b111111101100011010001;
		14'b00101010101110:	sigmoid = 21'b111111101100011100100;
		14'b00101010101111:	sigmoid = 21'b111111101100011111000;
		14'b00101010110000:	sigmoid = 21'b111111101100100001011;
		14'b00101010110001:	sigmoid = 21'b111111101100100011110;
		14'b00101010110010:	sigmoid = 21'b111111101100100110010;
		14'b00101010110011:	sigmoid = 21'b111111101100101000101;
		14'b00101010110100:	sigmoid = 21'b111111101100101011000;
		14'b00101010110101:	sigmoid = 21'b111111101100101101100;
		14'b00101010110110:	sigmoid = 21'b111111101100101111111;
		14'b00101010110111:	sigmoid = 21'b111111101100110010010;
		14'b00101010111000:	sigmoid = 21'b111111101100110100101;
		14'b00101010111001:	sigmoid = 21'b111111101100110111000;
		14'b00101010111010:	sigmoid = 21'b111111101100111001011;
		14'b00101010111011:	sigmoid = 21'b111111101100111011110;
		14'b00101010111100:	sigmoid = 21'b111111101100111110001;
		14'b00101010111101:	sigmoid = 21'b111111101101000000100;
		14'b00101010111110:	sigmoid = 21'b111111101101000010111;
		14'b00101010111111:	sigmoid = 21'b111111101101000101010;
		14'b00101011000000:	sigmoid = 21'b111111101101000111101;
		14'b00101011000001:	sigmoid = 21'b111111101101001001111;
		14'b00101011000010:	sigmoid = 21'b111111101101001100010;
		14'b00101011000011:	sigmoid = 21'b111111101101001110101;
		14'b00101011000100:	sigmoid = 21'b111111101101010000111;
		14'b00101011000101:	sigmoid = 21'b111111101101010011010;
		14'b00101011000110:	sigmoid = 21'b111111101101010101101;
		14'b00101011000111:	sigmoid = 21'b111111101101010111111;
		14'b00101011001000:	sigmoid = 21'b111111101101011010010;
		14'b00101011001001:	sigmoid = 21'b111111101101011100100;
		14'b00101011001010:	sigmoid = 21'b111111101101011110111;
		14'b00101011001011:	sigmoid = 21'b111111101101100001001;
		14'b00101011001100:	sigmoid = 21'b111111101101100011011;
		14'b00101011001101:	sigmoid = 21'b111111101101100101110;
		14'b00101011001110:	sigmoid = 21'b111111101101101000000;
		14'b00101011001111:	sigmoid = 21'b111111101101101010010;
		14'b00101011010000:	sigmoid = 21'b111111101101101100101;
		14'b00101011010001:	sigmoid = 21'b111111101101101110111;
		14'b00101011010010:	sigmoid = 21'b111111101101110001001;
		14'b00101011010011:	sigmoid = 21'b111111101101110011011;
		14'b00101011010100:	sigmoid = 21'b111111101101110101101;
		14'b00101011010101:	sigmoid = 21'b111111101101110111111;
		14'b00101011010110:	sigmoid = 21'b111111101101111010001;
		14'b00101011010111:	sigmoid = 21'b111111101101111100011;
		14'b00101011011000:	sigmoid = 21'b111111101101111110101;
		14'b00101011011001:	sigmoid = 21'b111111101110000000111;
		14'b00101011011010:	sigmoid = 21'b111111101110000011001;
		14'b00101011011011:	sigmoid = 21'b111111101110000101011;
		14'b00101011011100:	sigmoid = 21'b111111101110000111101;
		14'b00101011011101:	sigmoid = 21'b111111101110001001111;
		14'b00101011011110:	sigmoid = 21'b111111101110001100000;
		14'b00101011011111:	sigmoid = 21'b111111101110001110010;
		14'b00101011100000:	sigmoid = 21'b111111101110010000100;
		14'b00101011100001:	sigmoid = 21'b111111101110010010101;
		14'b00101011100010:	sigmoid = 21'b111111101110010100111;
		14'b00101011100011:	sigmoid = 21'b111111101110010111001;
		14'b00101011100100:	sigmoid = 21'b111111101110011001010;
		14'b00101011100101:	sigmoid = 21'b111111101110011011100;
		14'b00101011100110:	sigmoid = 21'b111111101110011101101;
		14'b00101011100111:	sigmoid = 21'b111111101110011111111;
		14'b00101011101000:	sigmoid = 21'b111111101110100010000;
		14'b00101011101001:	sigmoid = 21'b111111101110100100001;
		14'b00101011101010:	sigmoid = 21'b111111101110100110011;
		14'b00101011101011:	sigmoid = 21'b111111101110101000100;
		14'b00101011101100:	sigmoid = 21'b111111101110101010101;
		14'b00101011101101:	sigmoid = 21'b111111101110101100110;
		14'b00101011101110:	sigmoid = 21'b111111101110101111000;
		14'b00101011101111:	sigmoid = 21'b111111101110110001001;
		14'b00101011110000:	sigmoid = 21'b111111101110110011010;
		14'b00101011110001:	sigmoid = 21'b111111101110110101011;
		14'b00101011110010:	sigmoid = 21'b111111101110110111100;
		14'b00101011110011:	sigmoid = 21'b111111101110111001101;
		14'b00101011110100:	sigmoid = 21'b111111101110111011110;
		14'b00101011110101:	sigmoid = 21'b111111101110111101111;
		14'b00101011110110:	sigmoid = 21'b111111101111000000000;
		14'b00101011110111:	sigmoid = 21'b111111101111000010001;
		14'b00101011111000:	sigmoid = 21'b111111101111000100010;
		14'b00101011111001:	sigmoid = 21'b111111101111000110011;
		14'b00101011111010:	sigmoid = 21'b111111101111001000100;
		14'b00101011111011:	sigmoid = 21'b111111101111001010100;
		14'b00101011111100:	sigmoid = 21'b111111101111001100101;
		14'b00101011111101:	sigmoid = 21'b111111101111001110110;
		14'b00101011111110:	sigmoid = 21'b111111101111010000111;
		14'b00101011111111:	sigmoid = 21'b111111101111010010111;
		14'b00101100000000:	sigmoid = 21'b111111101111010101000;
		14'b00101100000001:	sigmoid = 21'b111111101111010111000;
		14'b00101100000010:	sigmoid = 21'b111111101111011001001;
		14'b00101100000011:	sigmoid = 21'b111111101111011011001;
		14'b00101100000100:	sigmoid = 21'b111111101111011101010;
		14'b00101100000101:	sigmoid = 21'b111111101111011111010;
		14'b00101100000110:	sigmoid = 21'b111111101111100001011;
		14'b00101100000111:	sigmoid = 21'b111111101111100011011;
		14'b00101100001000:	sigmoid = 21'b111111101111100101100;
		14'b00101100001001:	sigmoid = 21'b111111101111100111100;
		14'b00101100001010:	sigmoid = 21'b111111101111101001100;
		14'b00101100001011:	sigmoid = 21'b111111101111101011101;
		14'b00101100001100:	sigmoid = 21'b111111101111101101101;
		14'b00101100001101:	sigmoid = 21'b111111101111101111101;
		14'b00101100001110:	sigmoid = 21'b111111101111110001101;
		14'b00101100001111:	sigmoid = 21'b111111101111110011101;
		14'b00101100010000:	sigmoid = 21'b111111101111110101101;
		14'b00101100010001:	sigmoid = 21'b111111101111110111101;
		14'b00101100010010:	sigmoid = 21'b111111101111111001110;
		14'b00101100010011:	sigmoid = 21'b111111101111111011110;
		14'b00101100010100:	sigmoid = 21'b111111101111111101110;
		14'b00101100010101:	sigmoid = 21'b111111101111111111101;
		14'b00101100010110:	sigmoid = 21'b111111110000000001101;
		14'b00101100010111:	sigmoid = 21'b111111110000000011101;
		14'b00101100011000:	sigmoid = 21'b111111110000000101101;
		14'b00101100011001:	sigmoid = 21'b111111110000000111101;
		14'b00101100011010:	sigmoid = 21'b111111110000001001101;
		14'b00101100011011:	sigmoid = 21'b111111110000001011101;
		14'b00101100011100:	sigmoid = 21'b111111110000001101100;
		14'b00101100011101:	sigmoid = 21'b111111110000001111100;
		14'b00101100011110:	sigmoid = 21'b111111110000010001100;
		14'b00101100011111:	sigmoid = 21'b111111110000010011011;
		14'b00101100100000:	sigmoid = 21'b111111110000010101011;
		14'b00101100100001:	sigmoid = 21'b111111110000010111011;
		14'b00101100100010:	sigmoid = 21'b111111110000011001010;
		14'b00101100100011:	sigmoid = 21'b111111110000011011010;
		14'b00101100100100:	sigmoid = 21'b111111110000011101001;
		14'b00101100100101:	sigmoid = 21'b111111110000011111001;
		14'b00101100100110:	sigmoid = 21'b111111110000100001000;
		14'b00101100100111:	sigmoid = 21'b111111110000100010111;
		14'b00101100101000:	sigmoid = 21'b111111110000100100111;
		14'b00101100101001:	sigmoid = 21'b111111110000100110110;
		14'b00101100101010:	sigmoid = 21'b111111110000101000110;
		14'b00101100101011:	sigmoid = 21'b111111110000101010101;
		14'b00101100101100:	sigmoid = 21'b111111110000101100100;
		14'b00101100101101:	sigmoid = 21'b111111110000101110011;
		14'b00101100101110:	sigmoid = 21'b111111110000110000011;
		14'b00101100101111:	sigmoid = 21'b111111110000110010010;
		14'b00101100110000:	sigmoid = 21'b111111110000110100001;
		14'b00101100110001:	sigmoid = 21'b111111110000110110000;
		14'b00101100110010:	sigmoid = 21'b111111110000110111111;
		14'b00101100110011:	sigmoid = 21'b111111110000111001110;
		14'b00101100110100:	sigmoid = 21'b111111110000111011101;
		14'b00101100110101:	sigmoid = 21'b111111110000111101100;
		14'b00101100110110:	sigmoid = 21'b111111110000111111011;
		14'b00101100110111:	sigmoid = 21'b111111110001000001010;
		14'b00101100111000:	sigmoid = 21'b111111110001000011001;
		14'b00101100111001:	sigmoid = 21'b111111110001000101000;
		14'b00101100111010:	sigmoid = 21'b111111110001000110111;
		14'b00101100111011:	sigmoid = 21'b111111110001001000101;
		14'b00101100111100:	sigmoid = 21'b111111110001001010100;
		14'b00101100111101:	sigmoid = 21'b111111110001001100011;
		14'b00101100111110:	sigmoid = 21'b111111110001001110010;
		14'b00101100111111:	sigmoid = 21'b111111110001010000000;
		14'b00101101000000:	sigmoid = 21'b111111110001010001111;
		14'b00101101000001:	sigmoid = 21'b111111110001010011110;
		14'b00101101000010:	sigmoid = 21'b111111110001010101100;
		14'b00101101000011:	sigmoid = 21'b111111110001010111011;
		14'b00101101000100:	sigmoid = 21'b111111110001011001010;
		14'b00101101000101:	sigmoid = 21'b111111110001011011000;
		14'b00101101000110:	sigmoid = 21'b111111110001011100111;
		14'b00101101000111:	sigmoid = 21'b111111110001011110101;
		14'b00101101001000:	sigmoid = 21'b111111110001100000100;
		14'b00101101001001:	sigmoid = 21'b111111110001100010010;
		14'b00101101001010:	sigmoid = 21'b111111110001100100000;
		14'b00101101001011:	sigmoid = 21'b111111110001100101111;
		14'b00101101001100:	sigmoid = 21'b111111110001100111101;
		14'b00101101001101:	sigmoid = 21'b111111110001101001011;
		14'b00101101001110:	sigmoid = 21'b111111110001101011010;
		14'b00101101001111:	sigmoid = 21'b111111110001101101000;
		14'b00101101010000:	sigmoid = 21'b111111110001101110110;
		14'b00101101010001:	sigmoid = 21'b111111110001110000100;
		14'b00101101010010:	sigmoid = 21'b111111110001110010011;
		14'b00101101010011:	sigmoid = 21'b111111110001110100001;
		14'b00101101010100:	sigmoid = 21'b111111110001110101111;
		14'b00101101010101:	sigmoid = 21'b111111110001110111101;
		14'b00101101010110:	sigmoid = 21'b111111110001111001011;
		14'b00101101010111:	sigmoid = 21'b111111110001111011001;
		14'b00101101011000:	sigmoid = 21'b111111110001111100111;
		14'b00101101011001:	sigmoid = 21'b111111110001111110101;
		14'b00101101011010:	sigmoid = 21'b111111110010000000011;
		14'b00101101011011:	sigmoid = 21'b111111110010000010001;
		14'b00101101011100:	sigmoid = 21'b111111110010000011111;
		14'b00101101011101:	sigmoid = 21'b111111110010000101101;
		14'b00101101011110:	sigmoid = 21'b111111110010000111011;
		14'b00101101011111:	sigmoid = 21'b111111110010001001000;
		14'b00101101100000:	sigmoid = 21'b111111110010001010110;
		14'b00101101100001:	sigmoid = 21'b111111110010001100100;
		14'b00101101100010:	sigmoid = 21'b111111110010001110010;
		14'b00101101100011:	sigmoid = 21'b111111110010001111111;
		14'b00101101100100:	sigmoid = 21'b111111110010010001101;
		14'b00101101100101:	sigmoid = 21'b111111110010010011011;
		14'b00101101100110:	sigmoid = 21'b111111110010010101000;
		14'b00101101100111:	sigmoid = 21'b111111110010010110110;
		14'b00101101101000:	sigmoid = 21'b111111110010011000100;
		14'b00101101101001:	sigmoid = 21'b111111110010011010001;
		14'b00101101101010:	sigmoid = 21'b111111110010011011111;
		14'b00101101101011:	sigmoid = 21'b111111110010011101100;
		14'b00101101101100:	sigmoid = 21'b111111110010011111010;
		14'b00101101101101:	sigmoid = 21'b111111110010100000111;
		14'b00101101101110:	sigmoid = 21'b111111110010100010101;
		14'b00101101101111:	sigmoid = 21'b111111110010100100010;
		14'b00101101110000:	sigmoid = 21'b111111110010100101111;
		14'b00101101110001:	sigmoid = 21'b111111110010100111101;
		14'b00101101110010:	sigmoid = 21'b111111110010101001010;
		14'b00101101110011:	sigmoid = 21'b111111110010101010111;
		14'b00101101110100:	sigmoid = 21'b111111110010101100101;
		14'b00101101110101:	sigmoid = 21'b111111110010101110010;
		14'b00101101110110:	sigmoid = 21'b111111110010101111111;
		14'b00101101110111:	sigmoid = 21'b111111110010110001100;
		14'b00101101111000:	sigmoid = 21'b111111110010110011001;
		14'b00101101111001:	sigmoid = 21'b111111110010110100111;
		14'b00101101111010:	sigmoid = 21'b111111110010110110100;
		14'b00101101111011:	sigmoid = 21'b111111110010111000001;
		14'b00101101111100:	sigmoid = 21'b111111110010111001110;
		14'b00101101111101:	sigmoid = 21'b111111110010111011011;
		14'b00101101111110:	sigmoid = 21'b111111110010111101000;
		14'b00101101111111:	sigmoid = 21'b111111110010111110101;
		14'b00101110000000:	sigmoid = 21'b111111110011000000010;
		14'b00101110000001:	sigmoid = 21'b111111110011000001111;
		14'b00101110000010:	sigmoid = 21'b111111110011000011100;
		14'b00101110000011:	sigmoid = 21'b111111110011000101001;
		14'b00101110000100:	sigmoid = 21'b111111110011000110110;
		14'b00101110000101:	sigmoid = 21'b111111110011001000010;
		14'b00101110000110:	sigmoid = 21'b111111110011001001111;
		14'b00101110000111:	sigmoid = 21'b111111110011001011100;
		14'b00101110001000:	sigmoid = 21'b111111110011001101001;
		14'b00101110001001:	sigmoid = 21'b111111110011001110101;
		14'b00101110001010:	sigmoid = 21'b111111110011010000010;
		14'b00101110001011:	sigmoid = 21'b111111110011010001111;
		14'b00101110001100:	sigmoid = 21'b111111110011010011100;
		14'b00101110001101:	sigmoid = 21'b111111110011010101000;
		14'b00101110001110:	sigmoid = 21'b111111110011010110101;
		14'b00101110001111:	sigmoid = 21'b111111110011011000001;
		14'b00101110010000:	sigmoid = 21'b111111110011011001110;
		14'b00101110010001:	sigmoid = 21'b111111110011011011011;
		14'b00101110010010:	sigmoid = 21'b111111110011011100111;
		14'b00101110010011:	sigmoid = 21'b111111110011011110100;
		14'b00101110010100:	sigmoid = 21'b111111110011100000000;
		14'b00101110010101:	sigmoid = 21'b111111110011100001100;
		14'b00101110010110:	sigmoid = 21'b111111110011100011001;
		14'b00101110010111:	sigmoid = 21'b111111110011100100101;
		14'b00101110011000:	sigmoid = 21'b111111110011100110010;
		14'b00101110011001:	sigmoid = 21'b111111110011100111110;
		14'b00101110011010:	sigmoid = 21'b111111110011101001010;
		14'b00101110011011:	sigmoid = 21'b111111110011101010111;
		14'b00101110011100:	sigmoid = 21'b111111110011101100011;
		14'b00101110011101:	sigmoid = 21'b111111110011101101111;
		14'b00101110011110:	sigmoid = 21'b111111110011101111011;
		14'b00101110011111:	sigmoid = 21'b111111110011110001000;
		14'b00101110100000:	sigmoid = 21'b111111110011110010100;
		14'b00101110100001:	sigmoid = 21'b111111110011110100000;
		14'b00101110100010:	sigmoid = 21'b111111110011110101100;
		14'b00101110100011:	sigmoid = 21'b111111110011110111000;
		14'b00101110100100:	sigmoid = 21'b111111110011111000100;
		14'b00101110100101:	sigmoid = 21'b111111110011111010000;
		14'b00101110100110:	sigmoid = 21'b111111110011111011100;
		14'b00101110100111:	sigmoid = 21'b111111110011111101000;
		14'b00101110101000:	sigmoid = 21'b111111110011111110100;
		14'b00101110101001:	sigmoid = 21'b111111110100000000000;
		14'b00101110101010:	sigmoid = 21'b111111110100000001100;
		14'b00101110101011:	sigmoid = 21'b111111110100000011000;
		14'b00101110101100:	sigmoid = 21'b111111110100000100100;
		14'b00101110101101:	sigmoid = 21'b111111110100000110000;
		14'b00101110101110:	sigmoid = 21'b111111110100000111100;
		14'b00101110101111:	sigmoid = 21'b111111110100001001000;
		14'b00101110110000:	sigmoid = 21'b111111110100001010100;
		14'b00101110110001:	sigmoid = 21'b111111110100001011111;
		14'b00101110110010:	sigmoid = 21'b111111110100001101011;
		14'b00101110110011:	sigmoid = 21'b111111110100001110111;
		14'b00101110110100:	sigmoid = 21'b111111110100010000011;
		14'b00101110110101:	sigmoid = 21'b111111110100010001110;
		14'b00101110110110:	sigmoid = 21'b111111110100010011010;
		14'b00101110110111:	sigmoid = 21'b111111110100010100110;
		14'b00101110111000:	sigmoid = 21'b111111110100010110001;
		14'b00101110111001:	sigmoid = 21'b111111110100010111101;
		14'b00101110111010:	sigmoid = 21'b111111110100011001000;
		14'b00101110111011:	sigmoid = 21'b111111110100011010100;
		14'b00101110111100:	sigmoid = 21'b111111110100011100000;
		14'b00101110111101:	sigmoid = 21'b111111110100011101011;
		14'b00101110111110:	sigmoid = 21'b111111110100011110111;
		14'b00101110111111:	sigmoid = 21'b111111110100100000010;
		14'b00101111000000:	sigmoid = 21'b111111110100100001110;
		14'b00101111000001:	sigmoid = 21'b111111110100100011001;
		14'b00101111000010:	sigmoid = 21'b111111110100100100100;
		14'b00101111000011:	sigmoid = 21'b111111110100100110000;
		14'b00101111000100:	sigmoid = 21'b111111110100100111011;
		14'b00101111000101:	sigmoid = 21'b111111110100101000110;
		14'b00101111000110:	sigmoid = 21'b111111110100101010010;
		14'b00101111000111:	sigmoid = 21'b111111110100101011101;
		14'b00101111001000:	sigmoid = 21'b111111110100101101000;
		14'b00101111001001:	sigmoid = 21'b111111110100101110100;
		14'b00101111001010:	sigmoid = 21'b111111110100101111111;
		14'b00101111001011:	sigmoid = 21'b111111110100110001010;
		14'b00101111001100:	sigmoid = 21'b111111110100110010101;
		14'b00101111001101:	sigmoid = 21'b111111110100110100000;
		14'b00101111001110:	sigmoid = 21'b111111110100110101100;
		14'b00101111001111:	sigmoid = 21'b111111110100110110111;
		14'b00101111010000:	sigmoid = 21'b111111110100111000010;
		14'b00101111010001:	sigmoid = 21'b111111110100111001101;
		14'b00101111010010:	sigmoid = 21'b111111110100111011000;
		14'b00101111010011:	sigmoid = 21'b111111110100111100011;
		14'b00101111010100:	sigmoid = 21'b111111110100111101110;
		14'b00101111010101:	sigmoid = 21'b111111110100111111001;
		14'b00101111010110:	sigmoid = 21'b111111110101000000100;
		14'b00101111010111:	sigmoid = 21'b111111110101000001111;
		14'b00101111011000:	sigmoid = 21'b111111110101000011010;
		14'b00101111011001:	sigmoid = 21'b111111110101000100101;
		14'b00101111011010:	sigmoid = 21'b111111110101000110000;
		14'b00101111011011:	sigmoid = 21'b111111110101000111010;
		14'b00101111011100:	sigmoid = 21'b111111110101001000101;
		14'b00101111011101:	sigmoid = 21'b111111110101001010000;
		14'b00101111011110:	sigmoid = 21'b111111110101001011011;
		14'b00101111011111:	sigmoid = 21'b111111110101001100110;
		14'b00101111100000:	sigmoid = 21'b111111110101001110000;
		14'b00101111100001:	sigmoid = 21'b111111110101001111011;
		14'b00101111100010:	sigmoid = 21'b111111110101010000110;
		14'b00101111100011:	sigmoid = 21'b111111110101010010001;
		14'b00101111100100:	sigmoid = 21'b111111110101010011011;
		14'b00101111100101:	sigmoid = 21'b111111110101010100110;
		14'b00101111100110:	sigmoid = 21'b111111110101010110001;
		14'b00101111100111:	sigmoid = 21'b111111110101010111011;
		14'b00101111101000:	sigmoid = 21'b111111110101011000110;
		14'b00101111101001:	sigmoid = 21'b111111110101011010000;
		14'b00101111101010:	sigmoid = 21'b111111110101011011011;
		14'b00101111101011:	sigmoid = 21'b111111110101011100101;
		14'b00101111101100:	sigmoid = 21'b111111110101011110000;
		14'b00101111101101:	sigmoid = 21'b111111110101011111010;
		14'b00101111101110:	sigmoid = 21'b111111110101100000101;
		14'b00101111101111:	sigmoid = 21'b111111110101100001111;
		14'b00101111110000:	sigmoid = 21'b111111110101100011010;
		14'b00101111110001:	sigmoid = 21'b111111110101100100100;
		14'b00101111110010:	sigmoid = 21'b111111110101100101111;
		14'b00101111110011:	sigmoid = 21'b111111110101100111001;
		14'b00101111110100:	sigmoid = 21'b111111110101101000011;
		14'b00101111110101:	sigmoid = 21'b111111110101101001110;
		14'b00101111110110:	sigmoid = 21'b111111110101101011000;
		14'b00101111110111:	sigmoid = 21'b111111110101101100010;
		14'b00101111111000:	sigmoid = 21'b111111110101101101101;
		14'b00101111111001:	sigmoid = 21'b111111110101101110111;
		14'b00101111111010:	sigmoid = 21'b111111110101110000001;
		14'b00101111111011:	sigmoid = 21'b111111110101110001011;
		14'b00101111111100:	sigmoid = 21'b111111110101110010101;
		14'b00101111111101:	sigmoid = 21'b111111110101110100000;
		14'b00101111111110:	sigmoid = 21'b111111110101110101010;
		14'b00101111111111:	sigmoid = 21'b111111110101110110100;
		14'b00110000000000:	sigmoid = 21'b111111110101110111110;
		14'b00110000000001:	sigmoid = 21'b111111110101111001000;
		14'b00110000000010:	sigmoid = 21'b111111110101111010010;
		14'b00110000000011:	sigmoid = 21'b111111110101111011100;
		14'b00110000000100:	sigmoid = 21'b111111110101111100110;
		14'b00110000000101:	sigmoid = 21'b111111110101111110000;
		14'b00110000000110:	sigmoid = 21'b111111110101111111010;
		14'b00110000000111:	sigmoid = 21'b111111110110000000100;
		14'b00110000001000:	sigmoid = 21'b111111110110000001110;
		14'b00110000001001:	sigmoid = 21'b111111110110000011000;
		14'b00110000001010:	sigmoid = 21'b111111110110000100010;
		14'b00110000001011:	sigmoid = 21'b111111110110000101100;
		14'b00110000001100:	sigmoid = 21'b111111110110000110110;
		14'b00110000001101:	sigmoid = 21'b111111110110001000000;
		14'b00110000001110:	sigmoid = 21'b111111110110001001010;
		14'b00110000001111:	sigmoid = 21'b111111110110001010011;
		14'b00110000010000:	sigmoid = 21'b111111110110001011101;
		14'b00110000010001:	sigmoid = 21'b111111110110001100111;
		14'b00110000010010:	sigmoid = 21'b111111110110001110001;
		14'b00110000010011:	sigmoid = 21'b111111110110001111010;
		14'b00110000010100:	sigmoid = 21'b111111110110010000100;
		14'b00110000010101:	sigmoid = 21'b111111110110010001110;
		14'b00110000010110:	sigmoid = 21'b111111110110010011000;
		14'b00110000010111:	sigmoid = 21'b111111110110010100001;
		14'b00110000011000:	sigmoid = 21'b111111110110010101011;
		14'b00110000011001:	sigmoid = 21'b111111110110010110101;
		14'b00110000011010:	sigmoid = 21'b111111110110010111110;
		14'b00110000011011:	sigmoid = 21'b111111110110011001000;
		14'b00110000011100:	sigmoid = 21'b111111110110011010001;
		14'b00110000011101:	sigmoid = 21'b111111110110011011011;
		14'b00110000011110:	sigmoid = 21'b111111110110011100100;
		14'b00110000011111:	sigmoid = 21'b111111110110011101110;
		14'b00110000100000:	sigmoid = 21'b111111110110011110111;
		14'b00110000100001:	sigmoid = 21'b111111110110100000001;
		14'b00110000100010:	sigmoid = 21'b111111110110100001010;
		14'b00110000100011:	sigmoid = 21'b111111110110100010100;
		14'b00110000100100:	sigmoid = 21'b111111110110100011101;
		14'b00110000100101:	sigmoid = 21'b111111110110100100111;
		14'b00110000100110:	sigmoid = 21'b111111110110100110000;
		14'b00110000100111:	sigmoid = 21'b111111110110100111001;
		14'b00110000101000:	sigmoid = 21'b111111110110101000011;
		14'b00110000101001:	sigmoid = 21'b111111110110101001100;
		14'b00110000101010:	sigmoid = 21'b111111110110101010101;
		14'b00110000101011:	sigmoid = 21'b111111110110101011111;
		14'b00110000101100:	sigmoid = 21'b111111110110101101000;
		14'b00110000101101:	sigmoid = 21'b111111110110101110001;
		14'b00110000101110:	sigmoid = 21'b111111110110101111011;
		14'b00110000101111:	sigmoid = 21'b111111110110110000100;
		14'b00110000110000:	sigmoid = 21'b111111110110110001101;
		14'b00110000110001:	sigmoid = 21'b111111110110110010110;
		14'b00110000110010:	sigmoid = 21'b111111110110110011111;
		14'b00110000110011:	sigmoid = 21'b111111110110110101001;
		14'b00110000110100:	sigmoid = 21'b111111110110110110010;
		14'b00110000110101:	sigmoid = 21'b111111110110110111011;
		14'b00110000110110:	sigmoid = 21'b111111110110111000100;
		14'b00110000110111:	sigmoid = 21'b111111110110111001101;
		14'b00110000111000:	sigmoid = 21'b111111110110111010110;
		14'b00110000111001:	sigmoid = 21'b111111110110111011111;
		14'b00110000111010:	sigmoid = 21'b111111110110111101000;
		14'b00110000111011:	sigmoid = 21'b111111110110111110001;
		14'b00110000111100:	sigmoid = 21'b111111110110111111010;
		14'b00110000111101:	sigmoid = 21'b111111110111000000011;
		14'b00110000111110:	sigmoid = 21'b111111110111000001100;
		14'b00110000111111:	sigmoid = 21'b111111110111000010101;
		14'b00110001000000:	sigmoid = 21'b111111110111000011110;
		14'b00110001000001:	sigmoid = 21'b111111110111000100111;
		14'b00110001000010:	sigmoid = 21'b111111110111000110000;
		14'b00110001000011:	sigmoid = 21'b111111110111000111001;
		14'b00110001000100:	sigmoid = 21'b111111110111001000010;
		14'b00110001000101:	sigmoid = 21'b111111110111001001010;
		14'b00110001000110:	sigmoid = 21'b111111110111001010011;
		14'b00110001000111:	sigmoid = 21'b111111110111001011100;
		14'b00110001001000:	sigmoid = 21'b111111110111001100101;
		14'b00110001001001:	sigmoid = 21'b111111110111001101110;
		14'b00110001001010:	sigmoid = 21'b111111110111001110110;
		14'b00110001001011:	sigmoid = 21'b111111110111001111111;
		14'b00110001001100:	sigmoid = 21'b111111110111010001000;
		14'b00110001001101:	sigmoid = 21'b111111110111010010001;
		14'b00110001001110:	sigmoid = 21'b111111110111010011001;
		14'b00110001001111:	sigmoid = 21'b111111110111010100010;
		14'b00110001010000:	sigmoid = 21'b111111110111010101011;
		14'b00110001010001:	sigmoid = 21'b111111110111010110011;
		14'b00110001010010:	sigmoid = 21'b111111110111010111100;
		14'b00110001010011:	sigmoid = 21'b111111110111011000100;
		14'b00110001010100:	sigmoid = 21'b111111110111011001101;
		14'b00110001010101:	sigmoid = 21'b111111110111011010110;
		14'b00110001010110:	sigmoid = 21'b111111110111011011110;
		14'b00110001010111:	sigmoid = 21'b111111110111011100111;
		14'b00110001011000:	sigmoid = 21'b111111110111011101111;
		14'b00110001011001:	sigmoid = 21'b111111110111011111000;
		14'b00110001011010:	sigmoid = 21'b111111110111100000000;
		14'b00110001011011:	sigmoid = 21'b111111110111100001001;
		14'b00110001011100:	sigmoid = 21'b111111110111100010001;
		14'b00110001011101:	sigmoid = 21'b111111110111100011010;
		14'b00110001011110:	sigmoid = 21'b111111110111100100010;
		14'b00110001011111:	sigmoid = 21'b111111110111100101010;
		14'b00110001100000:	sigmoid = 21'b111111110111100110011;
		14'b00110001100001:	sigmoid = 21'b111111110111100111011;
		14'b00110001100010:	sigmoid = 21'b111111110111101000100;
		14'b00110001100011:	sigmoid = 21'b111111110111101001100;
		14'b00110001100100:	sigmoid = 21'b111111110111101010100;
		14'b00110001100101:	sigmoid = 21'b111111110111101011100;
		14'b00110001100110:	sigmoid = 21'b111111110111101100101;
		14'b00110001100111:	sigmoid = 21'b111111110111101101101;
		14'b00110001101000:	sigmoid = 21'b111111110111101110101;
		14'b00110001101001:	sigmoid = 21'b111111110111101111110;
		14'b00110001101010:	sigmoid = 21'b111111110111110000110;
		14'b00110001101011:	sigmoid = 21'b111111110111110001110;
		14'b00110001101100:	sigmoid = 21'b111111110111110010110;
		14'b00110001101101:	sigmoid = 21'b111111110111110011110;
		14'b00110001101110:	sigmoid = 21'b111111110111110100111;
		14'b00110001101111:	sigmoid = 21'b111111110111110101111;
		14'b00110001110000:	sigmoid = 21'b111111110111110110111;
		14'b00110001110001:	sigmoid = 21'b111111110111110111111;
		14'b00110001110010:	sigmoid = 21'b111111110111111000111;
		14'b00110001110011:	sigmoid = 21'b111111110111111001111;
		14'b00110001110100:	sigmoid = 21'b111111110111111010111;
		14'b00110001110101:	sigmoid = 21'b111111110111111011111;
		14'b00110001110110:	sigmoid = 21'b111111110111111100111;
		14'b00110001110111:	sigmoid = 21'b111111110111111101111;
		14'b00110001111000:	sigmoid = 21'b111111110111111110111;
		14'b00110001111001:	sigmoid = 21'b111111110111111111111;
		14'b00110001111010:	sigmoid = 21'b111111111000000000111;
		14'b00110001111011:	sigmoid = 21'b111111111000000001111;
		14'b00110001111100:	sigmoid = 21'b111111111000000010111;
		14'b00110001111101:	sigmoid = 21'b111111111000000011111;
		14'b00110001111110:	sigmoid = 21'b111111111000000100111;
		14'b00110001111111:	sigmoid = 21'b111111111000000101111;
		14'b00110010000000:	sigmoid = 21'b111111111000000110111;
		14'b00110010000001:	sigmoid = 21'b111111111000000111111;
		14'b00110010000010:	sigmoid = 21'b111111111000001000111;
		14'b00110010000011:	sigmoid = 21'b111111111000001001110;
		14'b00110010000100:	sigmoid = 21'b111111111000001010110;
		14'b00110010000101:	sigmoid = 21'b111111111000001011110;
		14'b00110010000110:	sigmoid = 21'b111111111000001100110;
		14'b00110010000111:	sigmoid = 21'b111111111000001101110;
		14'b00110010001000:	sigmoid = 21'b111111111000001110101;
		14'b00110010001001:	sigmoid = 21'b111111111000001111101;
		14'b00110010001010:	sigmoid = 21'b111111111000010000101;
		14'b00110010001011:	sigmoid = 21'b111111111000010001101;
		14'b00110010001100:	sigmoid = 21'b111111111000010010100;
		14'b00110010001101:	sigmoid = 21'b111111111000010011100;
		14'b00110010001110:	sigmoid = 21'b111111111000010100100;
		14'b00110010001111:	sigmoid = 21'b111111111000010101011;
		14'b00110010010000:	sigmoid = 21'b111111111000010110011;
		14'b00110010010001:	sigmoid = 21'b111111111000010111011;
		14'b00110010010010:	sigmoid = 21'b111111111000011000010;
		14'b00110010010011:	sigmoid = 21'b111111111000011001010;
		14'b00110010010100:	sigmoid = 21'b111111111000011010001;
		14'b00110010010101:	sigmoid = 21'b111111111000011011001;
		14'b00110010010110:	sigmoid = 21'b111111111000011100000;
		14'b00110010010111:	sigmoid = 21'b111111111000011101000;
		14'b00110010011000:	sigmoid = 21'b111111111000011110000;
		14'b00110010011001:	sigmoid = 21'b111111111000011110111;
		14'b00110010011010:	sigmoid = 21'b111111111000011111111;
		14'b00110010011011:	sigmoid = 21'b111111111000100000110;
		14'b00110010011100:	sigmoid = 21'b111111111000100001101;
		14'b00110010011101:	sigmoid = 21'b111111111000100010101;
		14'b00110010011110:	sigmoid = 21'b111111111000100011100;
		14'b00110010011111:	sigmoid = 21'b111111111000100100100;
		14'b00110010100000:	sigmoid = 21'b111111111000100101011;
		14'b00110010100001:	sigmoid = 21'b111111111000100110011;
		14'b00110010100010:	sigmoid = 21'b111111111000100111010;
		14'b00110010100011:	sigmoid = 21'b111111111000101000001;
		14'b00110010100100:	sigmoid = 21'b111111111000101001001;
		14'b00110010100101:	sigmoid = 21'b111111111000101010000;
		14'b00110010100110:	sigmoid = 21'b111111111000101010111;
		14'b00110010100111:	sigmoid = 21'b111111111000101011111;
		14'b00110010101000:	sigmoid = 21'b111111111000101100110;
		14'b00110010101001:	sigmoid = 21'b111111111000101101101;
		14'b00110010101010:	sigmoid = 21'b111111111000101110101;
		14'b00110010101011:	sigmoid = 21'b111111111000101111100;
		14'b00110010101100:	sigmoid = 21'b111111111000110000011;
		14'b00110010101101:	sigmoid = 21'b111111111000110001010;
		14'b00110010101110:	sigmoid = 21'b111111111000110010001;
		14'b00110010101111:	sigmoid = 21'b111111111000110011001;
		14'b00110010110000:	sigmoid = 21'b111111111000110100000;
		14'b00110010110001:	sigmoid = 21'b111111111000110100111;
		14'b00110010110010:	sigmoid = 21'b111111111000110101110;
		14'b00110010110011:	sigmoid = 21'b111111111000110110101;
		14'b00110010110100:	sigmoid = 21'b111111111000110111100;
		14'b00110010110101:	sigmoid = 21'b111111111000111000100;
		14'b00110010110110:	sigmoid = 21'b111111111000111001011;
		14'b00110010110111:	sigmoid = 21'b111111111000111010010;
		14'b00110010111000:	sigmoid = 21'b111111111000111011001;
		14'b00110010111001:	sigmoid = 21'b111111111000111100000;
		14'b00110010111010:	sigmoid = 21'b111111111000111100111;
		14'b00110010111011:	sigmoid = 21'b111111111000111101110;
		14'b00110010111100:	sigmoid = 21'b111111111000111110101;
		14'b00110010111101:	sigmoid = 21'b111111111000111111100;
		14'b00110010111110:	sigmoid = 21'b111111111001000000011;
		14'b00110010111111:	sigmoid = 21'b111111111001000001010;
		14'b00110011000000:	sigmoid = 21'b111111111001000010001;
		14'b00110011000001:	sigmoid = 21'b111111111001000011000;
		14'b00110011000010:	sigmoid = 21'b111111111001000011111;
		14'b00110011000011:	sigmoid = 21'b111111111001000100110;
		14'b00110011000100:	sigmoid = 21'b111111111001000101101;
		14'b00110011000101:	sigmoid = 21'b111111111001000110011;
		14'b00110011000110:	sigmoid = 21'b111111111001000111010;
		14'b00110011000111:	sigmoid = 21'b111111111001001000001;
		14'b00110011001000:	sigmoid = 21'b111111111001001001000;
		14'b00110011001001:	sigmoid = 21'b111111111001001001111;
		14'b00110011001010:	sigmoid = 21'b111111111001001010110;
		14'b00110011001011:	sigmoid = 21'b111111111001001011101;
		14'b00110011001100:	sigmoid = 21'b111111111001001100011;
		14'b00110011001101:	sigmoid = 21'b111111111001001101010;
		14'b00110011001110:	sigmoid = 21'b111111111001001110001;
		14'b00110011001111:	sigmoid = 21'b111111111001001111000;
		14'b00110011010000:	sigmoid = 21'b111111111001001111110;
		14'b00110011010001:	sigmoid = 21'b111111111001010000101;
		14'b00110011010010:	sigmoid = 21'b111111111001010001100;
		14'b00110011010011:	sigmoid = 21'b111111111001010010011;
		14'b00110011010100:	sigmoid = 21'b111111111001010011001;
		14'b00110011010101:	sigmoid = 21'b111111111001010100000;
		14'b00110011010110:	sigmoid = 21'b111111111001010100111;
		14'b00110011010111:	sigmoid = 21'b111111111001010101101;
		14'b00110011011000:	sigmoid = 21'b111111111001010110100;
		14'b00110011011001:	sigmoid = 21'b111111111001010111011;
		14'b00110011011010:	sigmoid = 21'b111111111001011000001;
		14'b00110011011011:	sigmoid = 21'b111111111001011001000;
		14'b00110011011100:	sigmoid = 21'b111111111001011001110;
		14'b00110011011101:	sigmoid = 21'b111111111001011010101;
		14'b00110011011110:	sigmoid = 21'b111111111001011011011;
		14'b00110011011111:	sigmoid = 21'b111111111001011100010;
		14'b00110011100000:	sigmoid = 21'b111111111001011101001;
		14'b00110011100001:	sigmoid = 21'b111111111001011101111;
		14'b00110011100010:	sigmoid = 21'b111111111001011110110;
		14'b00110011100011:	sigmoid = 21'b111111111001011111100;
		14'b00110011100100:	sigmoid = 21'b111111111001100000011;
		14'b00110011100101:	sigmoid = 21'b111111111001100001001;
		14'b00110011100110:	sigmoid = 21'b111111111001100010000;
		14'b00110011100111:	sigmoid = 21'b111111111001100010110;
		14'b00110011101000:	sigmoid = 21'b111111111001100011100;
		14'b00110011101001:	sigmoid = 21'b111111111001100100011;
		14'b00110011101010:	sigmoid = 21'b111111111001100101001;
		14'b00110011101011:	sigmoid = 21'b111111111001100110000;
		14'b00110011101100:	sigmoid = 21'b111111111001100110110;
		14'b00110011101101:	sigmoid = 21'b111111111001100111100;
		14'b00110011101110:	sigmoid = 21'b111111111001101000011;
		14'b00110011101111:	sigmoid = 21'b111111111001101001001;
		14'b00110011110000:	sigmoid = 21'b111111111001101010000;
		14'b00110011110001:	sigmoid = 21'b111111111001101010110;
		14'b00110011110010:	sigmoid = 21'b111111111001101011100;
		14'b00110011110011:	sigmoid = 21'b111111111001101100010;
		14'b00110011110100:	sigmoid = 21'b111111111001101101001;
		14'b00110011110101:	sigmoid = 21'b111111111001101101111;
		14'b00110011110110:	sigmoid = 21'b111111111001101110101;
		14'b00110011110111:	sigmoid = 21'b111111111001101111100;
		14'b00110011111000:	sigmoid = 21'b111111111001110000010;
		14'b00110011111001:	sigmoid = 21'b111111111001110001000;
		14'b00110011111010:	sigmoid = 21'b111111111001110001110;
		14'b00110011111011:	sigmoid = 21'b111111111001110010100;
		14'b00110011111100:	sigmoid = 21'b111111111001110011011;
		14'b00110011111101:	sigmoid = 21'b111111111001110100001;
		14'b00110011111110:	sigmoid = 21'b111111111001110100111;
		14'b00110011111111:	sigmoid = 21'b111111111001110101101;
		14'b00110100000000:	sigmoid = 21'b111111111001110110011;
		14'b00110100000001:	sigmoid = 21'b111111111001110111001;
		14'b00110100000010:	sigmoid = 21'b111111111001111000000;
		14'b00110100000011:	sigmoid = 21'b111111111001111000110;
		14'b00110100000100:	sigmoid = 21'b111111111001111001100;
		14'b00110100000101:	sigmoid = 21'b111111111001111010010;
		14'b00110100000110:	sigmoid = 21'b111111111001111011000;
		14'b00110100000111:	sigmoid = 21'b111111111001111011110;
		14'b00110100001000:	sigmoid = 21'b111111111001111100100;
		14'b00110100001001:	sigmoid = 21'b111111111001111101010;
		14'b00110100001010:	sigmoid = 21'b111111111001111110000;
		14'b00110100001011:	sigmoid = 21'b111111111001111110110;
		14'b00110100001100:	sigmoid = 21'b111111111001111111100;
		14'b00110100001101:	sigmoid = 21'b111111111010000000010;
		14'b00110100001110:	sigmoid = 21'b111111111010000001000;
		14'b00110100001111:	sigmoid = 21'b111111111010000001110;
		14'b00110100010000:	sigmoid = 21'b111111111010000010100;
		14'b00110100010001:	sigmoid = 21'b111111111010000011010;
		14'b00110100010010:	sigmoid = 21'b111111111010000100000;
		14'b00110100010011:	sigmoid = 21'b111111111010000100110;
		14'b00110100010100:	sigmoid = 21'b111111111010000101100;
		14'b00110100010101:	sigmoid = 21'b111111111010000110010;
		14'b00110100010110:	sigmoid = 21'b111111111010000111000;
		14'b00110100010111:	sigmoid = 21'b111111111010000111101;
		14'b00110100011000:	sigmoid = 21'b111111111010001000011;
		14'b00110100011001:	sigmoid = 21'b111111111010001001001;
		14'b00110100011010:	sigmoid = 21'b111111111010001001111;
		14'b00110100011011:	sigmoid = 21'b111111111010001010101;
		14'b00110100011100:	sigmoid = 21'b111111111010001011011;
		14'b00110100011101:	sigmoid = 21'b111111111010001100000;
		14'b00110100011110:	sigmoid = 21'b111111111010001100110;
		14'b00110100011111:	sigmoid = 21'b111111111010001101100;
		14'b00110100100000:	sigmoid = 21'b111111111010001110010;
		14'b00110100100001:	sigmoid = 21'b111111111010001111000;
		14'b00110100100010:	sigmoid = 21'b111111111010001111101;
		14'b00110100100011:	sigmoid = 21'b111111111010010000011;
		14'b00110100100100:	sigmoid = 21'b111111111010010001001;
		14'b00110100100101:	sigmoid = 21'b111111111010010001110;
		14'b00110100100110:	sigmoid = 21'b111111111010010010100;
		14'b00110100100111:	sigmoid = 21'b111111111010010011010;
		14'b00110100101000:	sigmoid = 21'b111111111010010100000;
		14'b00110100101001:	sigmoid = 21'b111111111010010100101;
		14'b00110100101010:	sigmoid = 21'b111111111010010101011;
		14'b00110100101011:	sigmoid = 21'b111111111010010110001;
		14'b00110100101100:	sigmoid = 21'b111111111010010110110;
		14'b00110100101101:	sigmoid = 21'b111111111010010111100;
		14'b00110100101110:	sigmoid = 21'b111111111010011000001;
		14'b00110100101111:	sigmoid = 21'b111111111010011000111;
		14'b00110100110000:	sigmoid = 21'b111111111010011001101;
		14'b00110100110001:	sigmoid = 21'b111111111010011010010;
		14'b00110100110010:	sigmoid = 21'b111111111010011011000;
		14'b00110100110011:	sigmoid = 21'b111111111010011011101;
		14'b00110100110100:	sigmoid = 21'b111111111010011100011;
		14'b00110100110101:	sigmoid = 21'b111111111010011101000;
		14'b00110100110110:	sigmoid = 21'b111111111010011101110;
		14'b00110100110111:	sigmoid = 21'b111111111010011110100;
		14'b00110100111000:	sigmoid = 21'b111111111010011111001;
		14'b00110100111001:	sigmoid = 21'b111111111010011111111;
		14'b00110100111010:	sigmoid = 21'b111111111010100000100;
		14'b00110100111011:	sigmoid = 21'b111111111010100001001;
		14'b00110100111100:	sigmoid = 21'b111111111010100001111;
		14'b00110100111101:	sigmoid = 21'b111111111010100010100;
		14'b00110100111110:	sigmoid = 21'b111111111010100011010;
		14'b00110100111111:	sigmoid = 21'b111111111010100011111;
		14'b00110101000000:	sigmoid = 21'b111111111010100100101;
		14'b00110101000001:	sigmoid = 21'b111111111010100101010;
		14'b00110101000010:	sigmoid = 21'b111111111010100110000;
		14'b00110101000011:	sigmoid = 21'b111111111010100110101;
		14'b00110101000100:	sigmoid = 21'b111111111010100111010;
		14'b00110101000101:	sigmoid = 21'b111111111010101000000;
		14'b00110101000110:	sigmoid = 21'b111111111010101000101;
		14'b00110101000111:	sigmoid = 21'b111111111010101001010;
		14'b00110101001000:	sigmoid = 21'b111111111010101010000;
		14'b00110101001001:	sigmoid = 21'b111111111010101010101;
		14'b00110101001010:	sigmoid = 21'b111111111010101011010;
		14'b00110101001011:	sigmoid = 21'b111111111010101100000;
		14'b00110101001100:	sigmoid = 21'b111111111010101100101;
		14'b00110101001101:	sigmoid = 21'b111111111010101101010;
		14'b00110101001110:	sigmoid = 21'b111111111010101110000;
		14'b00110101001111:	sigmoid = 21'b111111111010101110101;
		14'b00110101010000:	sigmoid = 21'b111111111010101111010;
		14'b00110101010001:	sigmoid = 21'b111111111010101111111;
		14'b00110101010010:	sigmoid = 21'b111111111010110000101;
		14'b00110101010011:	sigmoid = 21'b111111111010110001010;
		14'b00110101010100:	sigmoid = 21'b111111111010110001111;
		14'b00110101010101:	sigmoid = 21'b111111111010110010100;
		14'b00110101010110:	sigmoid = 21'b111111111010110011001;
		14'b00110101010111:	sigmoid = 21'b111111111010110011111;
		14'b00110101011000:	sigmoid = 21'b111111111010110100100;
		14'b00110101011001:	sigmoid = 21'b111111111010110101001;
		14'b00110101011010:	sigmoid = 21'b111111111010110101110;
		14'b00110101011011:	sigmoid = 21'b111111111010110110011;
		14'b00110101011100:	sigmoid = 21'b111111111010110111000;
		14'b00110101011101:	sigmoid = 21'b111111111010110111110;
		14'b00110101011110:	sigmoid = 21'b111111111010111000011;
		14'b00110101011111:	sigmoid = 21'b111111111010111001000;
		14'b00110101100000:	sigmoid = 21'b111111111010111001101;
		14'b00110101100001:	sigmoid = 21'b111111111010111010010;
		14'b00110101100010:	sigmoid = 21'b111111111010111010111;
		14'b00110101100011:	sigmoid = 21'b111111111010111011100;
		14'b00110101100100:	sigmoid = 21'b111111111010111100001;
		14'b00110101100101:	sigmoid = 21'b111111111010111100110;
		14'b00110101100110:	sigmoid = 21'b111111111010111101011;
		14'b00110101100111:	sigmoid = 21'b111111111010111110000;
		14'b00110101101000:	sigmoid = 21'b111111111010111110101;
		14'b00110101101001:	sigmoid = 21'b111111111010111111010;
		14'b00110101101010:	sigmoid = 21'b111111111010111111111;
		14'b00110101101011:	sigmoid = 21'b111111111011000000100;
		14'b00110101101100:	sigmoid = 21'b111111111011000001001;
		14'b00110101101101:	sigmoid = 21'b111111111011000001110;
		14'b00110101101110:	sigmoid = 21'b111111111011000010011;
		14'b00110101101111:	sigmoid = 21'b111111111011000011000;
		14'b00110101110000:	sigmoid = 21'b111111111011000011101;
		14'b00110101110001:	sigmoid = 21'b111111111011000100010;
		14'b00110101110010:	sigmoid = 21'b111111111011000100111;
		14'b00110101110011:	sigmoid = 21'b111111111011000101100;
		14'b00110101110100:	sigmoid = 21'b111111111011000110001;
		14'b00110101110101:	sigmoid = 21'b111111111011000110110;
		14'b00110101110110:	sigmoid = 21'b111111111011000111011;
		14'b00110101110111:	sigmoid = 21'b111111111011000111111;
		14'b00110101111000:	sigmoid = 21'b111111111011001000100;
		14'b00110101111001:	sigmoid = 21'b111111111011001001001;
		14'b00110101111010:	sigmoid = 21'b111111111011001001110;
		14'b00110101111011:	sigmoid = 21'b111111111011001010011;
		14'b00110101111100:	sigmoid = 21'b111111111011001011000;
		14'b00110101111101:	sigmoid = 21'b111111111011001011100;
		14'b00110101111110:	sigmoid = 21'b111111111011001100001;
		14'b00110101111111:	sigmoid = 21'b111111111011001100110;
		14'b00110110000000:	sigmoid = 21'b111111111011001101011;
		14'b00110110000001:	sigmoid = 21'b111111111011001110000;
		14'b00110110000010:	sigmoid = 21'b111111111011001110100;
		14'b00110110000011:	sigmoid = 21'b111111111011001111001;
		14'b00110110000100:	sigmoid = 21'b111111111011001111110;
		14'b00110110000101:	sigmoid = 21'b111111111011010000011;
		14'b00110110000110:	sigmoid = 21'b111111111011010000111;
		14'b00110110000111:	sigmoid = 21'b111111111011010001100;
		14'b00110110001000:	sigmoid = 21'b111111111011010010001;
		14'b00110110001001:	sigmoid = 21'b111111111011010010110;
		14'b00110110001010:	sigmoid = 21'b111111111011010011010;
		14'b00110110001011:	sigmoid = 21'b111111111011010011111;
		14'b00110110001100:	sigmoid = 21'b111111111011010100100;
		14'b00110110001101:	sigmoid = 21'b111111111011010101000;
		14'b00110110001110:	sigmoid = 21'b111111111011010101101;
		14'b00110110001111:	sigmoid = 21'b111111111011010110010;
		14'b00110110010000:	sigmoid = 21'b111111111011010110110;
		14'b00110110010001:	sigmoid = 21'b111111111011010111011;
		14'b00110110010010:	sigmoid = 21'b111111111011010111111;
		14'b00110110010011:	sigmoid = 21'b111111111011011000100;
		14'b00110110010100:	sigmoid = 21'b111111111011011001001;
		14'b00110110010101:	sigmoid = 21'b111111111011011001101;
		14'b00110110010110:	sigmoid = 21'b111111111011011010010;
		14'b00110110010111:	sigmoid = 21'b111111111011011010110;
		14'b00110110011000:	sigmoid = 21'b111111111011011011011;
		14'b00110110011001:	sigmoid = 21'b111111111011011100000;
		14'b00110110011010:	sigmoid = 21'b111111111011011100100;
		14'b00110110011011:	sigmoid = 21'b111111111011011101001;
		14'b00110110011100:	sigmoid = 21'b111111111011011101101;
		14'b00110110011101:	sigmoid = 21'b111111111011011110010;
		14'b00110110011110:	sigmoid = 21'b111111111011011110110;
		14'b00110110011111:	sigmoid = 21'b111111111011011111011;
		14'b00110110100000:	sigmoid = 21'b111111111011011111111;
		14'b00110110100001:	sigmoid = 21'b111111111011100000100;
		14'b00110110100010:	sigmoid = 21'b111111111011100001000;
		14'b00110110100011:	sigmoid = 21'b111111111011100001101;
		14'b00110110100100:	sigmoid = 21'b111111111011100010001;
		14'b00110110100101:	sigmoid = 21'b111111111011100010110;
		14'b00110110100110:	sigmoid = 21'b111111111011100011010;
		14'b00110110100111:	sigmoid = 21'b111111111011100011111;
		14'b00110110101000:	sigmoid = 21'b111111111011100100011;
		14'b00110110101001:	sigmoid = 21'b111111111011100100111;
		14'b00110110101010:	sigmoid = 21'b111111111011100101100;
		14'b00110110101011:	sigmoid = 21'b111111111011100110000;
		14'b00110110101100:	sigmoid = 21'b111111111011100110101;
		14'b00110110101101:	sigmoid = 21'b111111111011100111001;
		14'b00110110101110:	sigmoid = 21'b111111111011100111101;
		14'b00110110101111:	sigmoid = 21'b111111111011101000010;
		14'b00110110110000:	sigmoid = 21'b111111111011101000110;
		14'b00110110110001:	sigmoid = 21'b111111111011101001010;
		14'b00110110110010:	sigmoid = 21'b111111111011101001111;
		14'b00110110110011:	sigmoid = 21'b111111111011101010011;
		14'b00110110110100:	sigmoid = 21'b111111111011101010111;
		14'b00110110110101:	sigmoid = 21'b111111111011101011100;
		14'b00110110110110:	sigmoid = 21'b111111111011101100000;
		14'b00110110110111:	sigmoid = 21'b111111111011101100100;
		14'b00110110111000:	sigmoid = 21'b111111111011101101001;
		14'b00110110111001:	sigmoid = 21'b111111111011101101101;
		14'b00110110111010:	sigmoid = 21'b111111111011101110001;
		14'b00110110111011:	sigmoid = 21'b111111111011101110110;
		14'b00110110111100:	sigmoid = 21'b111111111011101111010;
		14'b00110110111101:	sigmoid = 21'b111111111011101111110;
		14'b00110110111110:	sigmoid = 21'b111111111011110000010;
		14'b00110110111111:	sigmoid = 21'b111111111011110000111;
		14'b00110111000000:	sigmoid = 21'b111111111011110001011;
		14'b00110111000001:	sigmoid = 21'b111111111011110001111;
		14'b00110111000010:	sigmoid = 21'b111111111011110010011;
		14'b00110111000011:	sigmoid = 21'b111111111011110010111;
		14'b00110111000100:	sigmoid = 21'b111111111011110011100;
		14'b00110111000101:	sigmoid = 21'b111111111011110100000;
		14'b00110111000110:	sigmoid = 21'b111111111011110100100;
		14'b00110111000111:	sigmoid = 21'b111111111011110101000;
		14'b00110111001000:	sigmoid = 21'b111111111011110101100;
		14'b00110111001001:	sigmoid = 21'b111111111011110110000;
		14'b00110111001010:	sigmoid = 21'b111111111011110110101;
		14'b00110111001011:	sigmoid = 21'b111111111011110111001;
		14'b00110111001100:	sigmoid = 21'b111111111011110111101;
		14'b00110111001101:	sigmoid = 21'b111111111011111000001;
		14'b00110111001110:	sigmoid = 21'b111111111011111000101;
		14'b00110111001111:	sigmoid = 21'b111111111011111001001;
		14'b00110111010000:	sigmoid = 21'b111111111011111001101;
		14'b00110111010001:	sigmoid = 21'b111111111011111010001;
		14'b00110111010010:	sigmoid = 21'b111111111011111010101;
		14'b00110111010011:	sigmoid = 21'b111111111011111011010;
		14'b00110111010100:	sigmoid = 21'b111111111011111011110;
		14'b00110111010101:	sigmoid = 21'b111111111011111100010;
		14'b00110111010110:	sigmoid = 21'b111111111011111100110;
		14'b00110111010111:	sigmoid = 21'b111111111011111101010;
		14'b00110111011000:	sigmoid = 21'b111111111011111101110;
		14'b00110111011001:	sigmoid = 21'b111111111011111110010;
		14'b00110111011010:	sigmoid = 21'b111111111011111110110;
		14'b00110111011011:	sigmoid = 21'b111111111011111111010;
		14'b00110111011100:	sigmoid = 21'b111111111011111111110;
		14'b00110111011101:	sigmoid = 21'b111111111100000000010;
		14'b00110111011110:	sigmoid = 21'b111111111100000000110;
		14'b00110111011111:	sigmoid = 21'b111111111100000001010;
		14'b00110111100000:	sigmoid = 21'b111111111100000001110;
		14'b00110111100001:	sigmoid = 21'b111111111100000010010;
		14'b00110111100010:	sigmoid = 21'b111111111100000010110;
		14'b00110111100011:	sigmoid = 21'b111111111100000011010;
		14'b00110111100100:	sigmoid = 21'b111111111100000011110;
		14'b00110111100101:	sigmoid = 21'b111111111100000100010;
		14'b00110111100110:	sigmoid = 21'b111111111100000100101;
		14'b00110111100111:	sigmoid = 21'b111111111100000101001;
		14'b00110111101000:	sigmoid = 21'b111111111100000101101;
		14'b00110111101001:	sigmoid = 21'b111111111100000110001;
		14'b00110111101010:	sigmoid = 21'b111111111100000110101;
		14'b00110111101011:	sigmoid = 21'b111111111100000111001;
		14'b00110111101100:	sigmoid = 21'b111111111100000111101;
		14'b00110111101101:	sigmoid = 21'b111111111100001000001;
		14'b00110111101110:	sigmoid = 21'b111111111100001000101;
		14'b00110111101111:	sigmoid = 21'b111111111100001001000;
		14'b00110111110000:	sigmoid = 21'b111111111100001001100;
		14'b00110111110001:	sigmoid = 21'b111111111100001010000;
		14'b00110111110010:	sigmoid = 21'b111111111100001010100;
		14'b00110111110011:	sigmoid = 21'b111111111100001011000;
		14'b00110111110100:	sigmoid = 21'b111111111100001011100;
		14'b00110111110101:	sigmoid = 21'b111111111100001011111;
		14'b00110111110110:	sigmoid = 21'b111111111100001100011;
		14'b00110111110111:	sigmoid = 21'b111111111100001100111;
		14'b00110111111000:	sigmoid = 21'b111111111100001101011;
		14'b00110111111001:	sigmoid = 21'b111111111100001101111;
		14'b00110111111010:	sigmoid = 21'b111111111100001110010;
		14'b00110111111011:	sigmoid = 21'b111111111100001110110;
		14'b00110111111100:	sigmoid = 21'b111111111100001111010;
		14'b00110111111101:	sigmoid = 21'b111111111100001111110;
		14'b00110111111110:	sigmoid = 21'b111111111100010000001;
		14'b00110111111111:	sigmoid = 21'b111111111100010000101;
		14'b00111000000000:	sigmoid = 21'b111111111100010001001;
		14'b00111000000001:	sigmoid = 21'b111111111100010001101;
		14'b00111000000010:	sigmoid = 21'b111111111100010010000;
		14'b00111000000011:	sigmoid = 21'b111111111100010010100;
		14'b00111000000100:	sigmoid = 21'b111111111100010011000;
		14'b00111000000101:	sigmoid = 21'b111111111100010011011;
		14'b00111000000110:	sigmoid = 21'b111111111100010011111;
		14'b00111000000111:	sigmoid = 21'b111111111100010100011;
		14'b00111000001000:	sigmoid = 21'b111111111100010100110;
		14'b00111000001001:	sigmoid = 21'b111111111100010101010;
		14'b00111000001010:	sigmoid = 21'b111111111100010101110;
		14'b00111000001011:	sigmoid = 21'b111111111100010110001;
		14'b00111000001100:	sigmoid = 21'b111111111100010110101;
		14'b00111000001101:	sigmoid = 21'b111111111100010111001;
		14'b00111000001110:	sigmoid = 21'b111111111100010111100;
		14'b00111000001111:	sigmoid = 21'b111111111100011000000;
		14'b00111000010000:	sigmoid = 21'b111111111100011000100;
		14'b00111000010001:	sigmoid = 21'b111111111100011000111;
		14'b00111000010010:	sigmoid = 21'b111111111100011001011;
		14'b00111000010011:	sigmoid = 21'b111111111100011001110;
		14'b00111000010100:	sigmoid = 21'b111111111100011010010;
		14'b00111000010101:	sigmoid = 21'b111111111100011010110;
		14'b00111000010110:	sigmoid = 21'b111111111100011011001;
		14'b00111000010111:	sigmoid = 21'b111111111100011011101;
		14'b00111000011000:	sigmoid = 21'b111111111100011100000;
		14'b00111000011001:	sigmoid = 21'b111111111100011100100;
		14'b00111000011010:	sigmoid = 21'b111111111100011100111;
		14'b00111000011011:	sigmoid = 21'b111111111100011101011;
		14'b00111000011100:	sigmoid = 21'b111111111100011101110;
		14'b00111000011101:	sigmoid = 21'b111111111100011110010;
		14'b00111000011110:	sigmoid = 21'b111111111100011110110;
		14'b00111000011111:	sigmoid = 21'b111111111100011111001;
		14'b00111000100000:	sigmoid = 21'b111111111100011111101;
		14'b00111000100001:	sigmoid = 21'b111111111100100000000;
		14'b00111000100010:	sigmoid = 21'b111111111100100000100;
		14'b00111000100011:	sigmoid = 21'b111111111100100000111;
		14'b00111000100100:	sigmoid = 21'b111111111100100001011;
		14'b00111000100101:	sigmoid = 21'b111111111100100001110;
		14'b00111000100110:	sigmoid = 21'b111111111100100010001;
		14'b00111000100111:	sigmoid = 21'b111111111100100010101;
		14'b00111000101000:	sigmoid = 21'b111111111100100011000;
		14'b00111000101001:	sigmoid = 21'b111111111100100011100;
		14'b00111000101010:	sigmoid = 21'b111111111100100011111;
		14'b00111000101011:	sigmoid = 21'b111111111100100100011;
		14'b00111000101100:	sigmoid = 21'b111111111100100100110;
		14'b00111000101101:	sigmoid = 21'b111111111100100101010;
		14'b00111000101110:	sigmoid = 21'b111111111100100101101;
		14'b00111000101111:	sigmoid = 21'b111111111100100110000;
		14'b00111000110000:	sigmoid = 21'b111111111100100110100;
		14'b00111000110001:	sigmoid = 21'b111111111100100110111;
		14'b00111000110010:	sigmoid = 21'b111111111100100111011;
		14'b00111000110011:	sigmoid = 21'b111111111100100111110;
		14'b00111000110100:	sigmoid = 21'b111111111100101000001;
		14'b00111000110101:	sigmoid = 21'b111111111100101000101;
		14'b00111000110110:	sigmoid = 21'b111111111100101001000;
		14'b00111000110111:	sigmoid = 21'b111111111100101001011;
		14'b00111000111000:	sigmoid = 21'b111111111100101001111;
		14'b00111000111001:	sigmoid = 21'b111111111100101010010;
		14'b00111000111010:	sigmoid = 21'b111111111100101010101;
		14'b00111000111011:	sigmoid = 21'b111111111100101011001;
		14'b00111000111100:	sigmoid = 21'b111111111100101011100;
		14'b00111000111101:	sigmoid = 21'b111111111100101011111;
		14'b00111000111110:	sigmoid = 21'b111111111100101100011;
		14'b00111000111111:	sigmoid = 21'b111111111100101100110;
		14'b00111001000000:	sigmoid = 21'b111111111100101101001;
		14'b00111001000001:	sigmoid = 21'b111111111100101101100;
		14'b00111001000010:	sigmoid = 21'b111111111100101110000;
		14'b00111001000011:	sigmoid = 21'b111111111100101110011;
		14'b00111001000100:	sigmoid = 21'b111111111100101110110;
		14'b00111001000101:	sigmoid = 21'b111111111100101111010;
		14'b00111001000110:	sigmoid = 21'b111111111100101111101;
		14'b00111001000111:	sigmoid = 21'b111111111100110000000;
		14'b00111001001000:	sigmoid = 21'b111111111100110000011;
		14'b00111001001001:	sigmoid = 21'b111111111100110000111;
		14'b00111001001010:	sigmoid = 21'b111111111100110001010;
		14'b00111001001011:	sigmoid = 21'b111111111100110001101;
		14'b00111001001100:	sigmoid = 21'b111111111100110010000;
		14'b00111001001101:	sigmoid = 21'b111111111100110010011;
		14'b00111001001110:	sigmoid = 21'b111111111100110010111;
		14'b00111001001111:	sigmoid = 21'b111111111100110011010;
		14'b00111001010000:	sigmoid = 21'b111111111100110011101;
		14'b00111001010001:	sigmoid = 21'b111111111100110100000;
		14'b00111001010010:	sigmoid = 21'b111111111100110100011;
		14'b00111001010011:	sigmoid = 21'b111111111100110100111;
		14'b00111001010100:	sigmoid = 21'b111111111100110101010;
		14'b00111001010101:	sigmoid = 21'b111111111100110101101;
		14'b00111001010110:	sigmoid = 21'b111111111100110110000;
		14'b00111001010111:	sigmoid = 21'b111111111100110110011;
		14'b00111001011000:	sigmoid = 21'b111111111100110110110;
		14'b00111001011001:	sigmoid = 21'b111111111100110111010;
		14'b00111001011010:	sigmoid = 21'b111111111100110111101;
		14'b00111001011011:	sigmoid = 21'b111111111100111000000;
		14'b00111001011100:	sigmoid = 21'b111111111100111000011;
		14'b00111001011101:	sigmoid = 21'b111111111100111000110;
		14'b00111001011110:	sigmoid = 21'b111111111100111001001;
		14'b00111001011111:	sigmoid = 21'b111111111100111001100;
		14'b00111001100000:	sigmoid = 21'b111111111100111001111;
		14'b00111001100001:	sigmoid = 21'b111111111100111010010;
		14'b00111001100010:	sigmoid = 21'b111111111100111010101;
		14'b00111001100011:	sigmoid = 21'b111111111100111011001;
		14'b00111001100100:	sigmoid = 21'b111111111100111011100;
		14'b00111001100101:	sigmoid = 21'b111111111100111011111;
		14'b00111001100110:	sigmoid = 21'b111111111100111100010;
		14'b00111001100111:	sigmoid = 21'b111111111100111100101;
		14'b00111001101000:	sigmoid = 21'b111111111100111101000;
		14'b00111001101001:	sigmoid = 21'b111111111100111101011;
		14'b00111001101010:	sigmoid = 21'b111111111100111101110;
		14'b00111001101011:	sigmoid = 21'b111111111100111110001;
		14'b00111001101100:	sigmoid = 21'b111111111100111110100;
		14'b00111001101101:	sigmoid = 21'b111111111100111110111;
		14'b00111001101110:	sigmoid = 21'b111111111100111111010;
		14'b00111001101111:	sigmoid = 21'b111111111100111111101;
		14'b00111001110000:	sigmoid = 21'b111111111101000000000;
		14'b00111001110001:	sigmoid = 21'b111111111101000000011;
		14'b00111001110010:	sigmoid = 21'b111111111101000000110;
		14'b00111001110011:	sigmoid = 21'b111111111101000001001;
		14'b00111001110100:	sigmoid = 21'b111111111101000001100;
		14'b00111001110101:	sigmoid = 21'b111111111101000001111;
		14'b00111001110110:	sigmoid = 21'b111111111101000010010;
		14'b00111001110111:	sigmoid = 21'b111111111101000010101;
		14'b00111001111000:	sigmoid = 21'b111111111101000011000;
		14'b00111001111001:	sigmoid = 21'b111111111101000011011;
		14'b00111001111010:	sigmoid = 21'b111111111101000011110;
		14'b00111001111011:	sigmoid = 21'b111111111101000100001;
		14'b00111001111100:	sigmoid = 21'b111111111101000100100;
		14'b00111001111101:	sigmoid = 21'b111111111101000100110;
		14'b00111001111110:	sigmoid = 21'b111111111101000101001;
		14'b00111001111111:	sigmoid = 21'b111111111101000101100;
		14'b00111010000000:	sigmoid = 21'b111111111101000101111;
		14'b00111010000001:	sigmoid = 21'b111111111101000110010;
		14'b00111010000010:	sigmoid = 21'b111111111101000110101;
		14'b00111010000011:	sigmoid = 21'b111111111101000111000;
		14'b00111010000100:	sigmoid = 21'b111111111101000111011;
		14'b00111010000101:	sigmoid = 21'b111111111101000111110;
		14'b00111010000110:	sigmoid = 21'b111111111101001000001;
		14'b00111010000111:	sigmoid = 21'b111111111101001000011;
		14'b00111010001000:	sigmoid = 21'b111111111101001000110;
		14'b00111010001001:	sigmoid = 21'b111111111101001001001;
		14'b00111010001010:	sigmoid = 21'b111111111101001001100;
		14'b00111010001011:	sigmoid = 21'b111111111101001001111;
		14'b00111010001100:	sigmoid = 21'b111111111101001010010;
		14'b00111010001101:	sigmoid = 21'b111111111101001010101;
		14'b00111010001110:	sigmoid = 21'b111111111101001010111;
		14'b00111010001111:	sigmoid = 21'b111111111101001011010;
		14'b00111010010000:	sigmoid = 21'b111111111101001011101;
		14'b00111010010001:	sigmoid = 21'b111111111101001100000;
		14'b00111010010010:	sigmoid = 21'b111111111101001100011;
		14'b00111010010011:	sigmoid = 21'b111111111101001100101;
		14'b00111010010100:	sigmoid = 21'b111111111101001101000;
		14'b00111010010101:	sigmoid = 21'b111111111101001101011;
		14'b00111010010110:	sigmoid = 21'b111111111101001101110;
		14'b00111010010111:	sigmoid = 21'b111111111101001110001;
		14'b00111010011000:	sigmoid = 21'b111111111101001110011;
		14'b00111010011001:	sigmoid = 21'b111111111101001110110;
		14'b00111010011010:	sigmoid = 21'b111111111101001111001;
		14'b00111010011011:	sigmoid = 21'b111111111101001111100;
		14'b00111010011100:	sigmoid = 21'b111111111101001111110;
		14'b00111010011101:	sigmoid = 21'b111111111101010000001;
		14'b00111010011110:	sigmoid = 21'b111111111101010000100;
		14'b00111010011111:	sigmoid = 21'b111111111101010000111;
		14'b00111010100000:	sigmoid = 21'b111111111101010001001;
		14'b00111010100001:	sigmoid = 21'b111111111101010001100;
		14'b00111010100010:	sigmoid = 21'b111111111101010001111;
		14'b00111010100011:	sigmoid = 21'b111111111101010010001;
		14'b00111010100100:	sigmoid = 21'b111111111101010010100;
		14'b00111010100101:	sigmoid = 21'b111111111101010010111;
		14'b00111010100110:	sigmoid = 21'b111111111101010011010;
		14'b00111010100111:	sigmoid = 21'b111111111101010011100;
		14'b00111010101000:	sigmoid = 21'b111111111101010011111;
		14'b00111010101001:	sigmoid = 21'b111111111101010100010;
		14'b00111010101010:	sigmoid = 21'b111111111101010100100;
		14'b00111010101011:	sigmoid = 21'b111111111101010100111;
		14'b00111010101100:	sigmoid = 21'b111111111101010101010;
		14'b00111010101101:	sigmoid = 21'b111111111101010101100;
		14'b00111010101110:	sigmoid = 21'b111111111101010101111;
		14'b00111010101111:	sigmoid = 21'b111111111101010110010;
		14'b00111010110000:	sigmoid = 21'b111111111101010110100;
		14'b00111010110001:	sigmoid = 21'b111111111101010110111;
		14'b00111010110010:	sigmoid = 21'b111111111101010111010;
		14'b00111010110011:	sigmoid = 21'b111111111101010111100;
		14'b00111010110100:	sigmoid = 21'b111111111101010111111;
		14'b00111010110101:	sigmoid = 21'b111111111101011000001;
		14'b00111010110110:	sigmoid = 21'b111111111101011000100;
		14'b00111010110111:	sigmoid = 21'b111111111101011000111;
		14'b00111010111000:	sigmoid = 21'b111111111101011001001;
		14'b00111010111001:	sigmoid = 21'b111111111101011001100;
		14'b00111010111010:	sigmoid = 21'b111111111101011001111;
		14'b00111010111011:	sigmoid = 21'b111111111101011010001;
		14'b00111010111100:	sigmoid = 21'b111111111101011010100;
		14'b00111010111101:	sigmoid = 21'b111111111101011010110;
		14'b00111010111110:	sigmoid = 21'b111111111101011011001;
		14'b00111010111111:	sigmoid = 21'b111111111101011011011;
		14'b00111011000000:	sigmoid = 21'b111111111101011011110;
		14'b00111011000001:	sigmoid = 21'b111111111101011100001;
		14'b00111011000010:	sigmoid = 21'b111111111101011100011;
		14'b00111011000011:	sigmoid = 21'b111111111101011100110;
		14'b00111011000100:	sigmoid = 21'b111111111101011101000;
		14'b00111011000101:	sigmoid = 21'b111111111101011101011;
		14'b00111011000110:	sigmoid = 21'b111111111101011101101;
		14'b00111011000111:	sigmoid = 21'b111111111101011110000;
		14'b00111011001000:	sigmoid = 21'b111111111101011110010;
		14'b00111011001001:	sigmoid = 21'b111111111101011110101;
		14'b00111011001010:	sigmoid = 21'b111111111101011110111;
		14'b00111011001011:	sigmoid = 21'b111111111101011111010;
		14'b00111011001100:	sigmoid = 21'b111111111101011111100;
		14'b00111011001101:	sigmoid = 21'b111111111101011111111;
		14'b00111011001110:	sigmoid = 21'b111111111101100000001;
		14'b00111011001111:	sigmoid = 21'b111111111101100000100;
		14'b00111011010000:	sigmoid = 21'b111111111101100000110;
		14'b00111011010001:	sigmoid = 21'b111111111101100001001;
		14'b00111011010010:	sigmoid = 21'b111111111101100001011;
		14'b00111011010011:	sigmoid = 21'b111111111101100001110;
		14'b00111011010100:	sigmoid = 21'b111111111101100010000;
		14'b00111011010101:	sigmoid = 21'b111111111101100010011;
		14'b00111011010110:	sigmoid = 21'b111111111101100010101;
		14'b00111011010111:	sigmoid = 21'b111111111101100011000;
		14'b00111011011000:	sigmoid = 21'b111111111101100011010;
		14'b00111011011001:	sigmoid = 21'b111111111101100011101;
		14'b00111011011010:	sigmoid = 21'b111111111101100011111;
		14'b00111011011011:	sigmoid = 21'b111111111101100100001;
		14'b00111011011100:	sigmoid = 21'b111111111101100100100;
		14'b00111011011101:	sigmoid = 21'b111111111101100100110;
		14'b00111011011110:	sigmoid = 21'b111111111101100101001;
		14'b00111011011111:	sigmoid = 21'b111111111101100101011;
		14'b00111011100000:	sigmoid = 21'b111111111101100101110;
		14'b00111011100001:	sigmoid = 21'b111111111101100110000;
		14'b00111011100010:	sigmoid = 21'b111111111101100110010;
		14'b00111011100011:	sigmoid = 21'b111111111101100110101;
		14'b00111011100100:	sigmoid = 21'b111111111101100110111;
		14'b00111011100101:	sigmoid = 21'b111111111101100111010;
		14'b00111011100110:	sigmoid = 21'b111111111101100111100;
		14'b00111011100111:	sigmoid = 21'b111111111101100111110;
		14'b00111011101000:	sigmoid = 21'b111111111101101000001;
		14'b00111011101001:	sigmoid = 21'b111111111101101000011;
		14'b00111011101010:	sigmoid = 21'b111111111101101000101;
		14'b00111011101011:	sigmoid = 21'b111111111101101001000;
		14'b00111011101100:	sigmoid = 21'b111111111101101001010;
		14'b00111011101101:	sigmoid = 21'b111111111101101001100;
		14'b00111011101110:	sigmoid = 21'b111111111101101001111;
		14'b00111011101111:	sigmoid = 21'b111111111101101010001;
		14'b00111011110000:	sigmoid = 21'b111111111101101010011;
		14'b00111011110001:	sigmoid = 21'b111111111101101010110;
		14'b00111011110010:	sigmoid = 21'b111111111101101011000;
		14'b00111011110011:	sigmoid = 21'b111111111101101011010;
		14'b00111011110100:	sigmoid = 21'b111111111101101011101;
		14'b00111011110101:	sigmoid = 21'b111111111101101011111;
		14'b00111011110110:	sigmoid = 21'b111111111101101100001;
		14'b00111011110111:	sigmoid = 21'b111111111101101100100;
		14'b00111011111000:	sigmoid = 21'b111111111101101100110;
		14'b00111011111001:	sigmoid = 21'b111111111101101101000;
		14'b00111011111010:	sigmoid = 21'b111111111101101101011;
		14'b00111011111011:	sigmoid = 21'b111111111101101101101;
		14'b00111011111100:	sigmoid = 21'b111111111101101101111;
		14'b00111011111101:	sigmoid = 21'b111111111101101110001;
		14'b00111011111110:	sigmoid = 21'b111111111101101110100;
		14'b00111011111111:	sigmoid = 21'b111111111101101110110;
		14'b00111100000000:	sigmoid = 21'b111111111101101111000;
		14'b00111100000001:	sigmoid = 21'b111111111101101111010;
		14'b00111100000010:	sigmoid = 21'b111111111101101111101;
		14'b00111100000011:	sigmoid = 21'b111111111101101111111;
		14'b00111100000100:	sigmoid = 21'b111111111101110000001;
		14'b00111100000101:	sigmoid = 21'b111111111101110000011;
		14'b00111100000110:	sigmoid = 21'b111111111101110000110;
		14'b00111100000111:	sigmoid = 21'b111111111101110001000;
		14'b00111100001000:	sigmoid = 21'b111111111101110001010;
		14'b00111100001001:	sigmoid = 21'b111111111101110001100;
		14'b00111100001010:	sigmoid = 21'b111111111101110001111;
		14'b00111100001011:	sigmoid = 21'b111111111101110010001;
		14'b00111100001100:	sigmoid = 21'b111111111101110010011;
		14'b00111100001101:	sigmoid = 21'b111111111101110010101;
		14'b00111100001110:	sigmoid = 21'b111111111101110010111;
		14'b00111100001111:	sigmoid = 21'b111111111101110011010;
		14'b00111100010000:	sigmoid = 21'b111111111101110011100;
		14'b00111100010001:	sigmoid = 21'b111111111101110011110;
		14'b00111100010010:	sigmoid = 21'b111111111101110100000;
		14'b00111100010011:	sigmoid = 21'b111111111101110100010;
		14'b00111100010100:	sigmoid = 21'b111111111101110100101;
		14'b00111100010101:	sigmoid = 21'b111111111101110100111;
		14'b00111100010110:	sigmoid = 21'b111111111101110101001;
		14'b00111100010111:	sigmoid = 21'b111111111101110101011;
		14'b00111100011000:	sigmoid = 21'b111111111101110101101;
		14'b00111100011001:	sigmoid = 21'b111111111101110101111;
		14'b00111100011010:	sigmoid = 21'b111111111101110110010;
		14'b00111100011011:	sigmoid = 21'b111111111101110110100;
		14'b00111100011100:	sigmoid = 21'b111111111101110110110;
		14'b00111100011101:	sigmoid = 21'b111111111101110111000;
		14'b00111100011110:	sigmoid = 21'b111111111101110111010;
		14'b00111100011111:	sigmoid = 21'b111111111101110111100;
		14'b00111100100000:	sigmoid = 21'b111111111101110111110;
		14'b00111100100001:	sigmoid = 21'b111111111101111000001;
		14'b00111100100010:	sigmoid = 21'b111111111101111000011;
		14'b00111100100011:	sigmoid = 21'b111111111101111000101;
		14'b00111100100100:	sigmoid = 21'b111111111101111000111;
		14'b00111100100101:	sigmoid = 21'b111111111101111001001;
		14'b00111100100110:	sigmoid = 21'b111111111101111001011;
		14'b00111100100111:	sigmoid = 21'b111111111101111001101;
		14'b00111100101000:	sigmoid = 21'b111111111101111001111;
		14'b00111100101001:	sigmoid = 21'b111111111101111010001;
		14'b00111100101010:	sigmoid = 21'b111111111101111010011;
		14'b00111100101011:	sigmoid = 21'b111111111101111010110;
		14'b00111100101100:	sigmoid = 21'b111111111101111011000;
		14'b00111100101101:	sigmoid = 21'b111111111101111011010;
		14'b00111100101110:	sigmoid = 21'b111111111101111011100;
		14'b00111100101111:	sigmoid = 21'b111111111101111011110;
		14'b00111100110000:	sigmoid = 21'b111111111101111100000;
		14'b00111100110001:	sigmoid = 21'b111111111101111100010;
		14'b00111100110010:	sigmoid = 21'b111111111101111100100;
		14'b00111100110011:	sigmoid = 21'b111111111101111100110;
		14'b00111100110100:	sigmoid = 21'b111111111101111101000;
		14'b00111100110101:	sigmoid = 21'b111111111101111101010;
		14'b00111100110110:	sigmoid = 21'b111111111101111101100;
		14'b00111100110111:	sigmoid = 21'b111111111101111101110;
		14'b00111100111000:	sigmoid = 21'b111111111101111110000;
		14'b00111100111001:	sigmoid = 21'b111111111101111110010;
		14'b00111100111010:	sigmoid = 21'b111111111101111110100;
		14'b00111100111011:	sigmoid = 21'b111111111101111110110;
		14'b00111100111100:	sigmoid = 21'b111111111101111111000;
		14'b00111100111101:	sigmoid = 21'b111111111101111111010;
		14'b00111100111110:	sigmoid = 21'b111111111101111111100;
		14'b00111100111111:	sigmoid = 21'b111111111101111111110;
		14'b00111101000000:	sigmoid = 21'b111111111110000000000;
		14'b00111101000001:	sigmoid = 21'b111111111110000000010;
		14'b00111101000010:	sigmoid = 21'b111111111110000000100;
		14'b00111101000011:	sigmoid = 21'b111111111110000000110;
		14'b00111101000100:	sigmoid = 21'b111111111110000001000;
		14'b00111101000101:	sigmoid = 21'b111111111110000001010;
		14'b00111101000110:	sigmoid = 21'b111111111110000001100;
		14'b00111101000111:	sigmoid = 21'b111111111110000001110;
		14'b00111101001000:	sigmoid = 21'b111111111110000010000;
		14'b00111101001001:	sigmoid = 21'b111111111110000010010;
		14'b00111101001010:	sigmoid = 21'b111111111110000010100;
		14'b00111101001011:	sigmoid = 21'b111111111110000010110;
		14'b00111101001100:	sigmoid = 21'b111111111110000011000;
		14'b00111101001101:	sigmoid = 21'b111111111110000011010;
		14'b00111101001110:	sigmoid = 21'b111111111110000011100;
		14'b00111101001111:	sigmoid = 21'b111111111110000011110;
		14'b00111101010000:	sigmoid = 21'b111111111110000100000;
		14'b00111101010001:	sigmoid = 21'b111111111110000100010;
		14'b00111101010010:	sigmoid = 21'b111111111110000100100;
		14'b00111101010011:	sigmoid = 21'b111111111110000100110;
		14'b00111101010100:	sigmoid = 21'b111111111110000101000;
		14'b00111101010101:	sigmoid = 21'b111111111110000101001;
		14'b00111101010110:	sigmoid = 21'b111111111110000101011;
		14'b00111101010111:	sigmoid = 21'b111111111110000101101;
		14'b00111101011000:	sigmoid = 21'b111111111110000101111;
		14'b00111101011001:	sigmoid = 21'b111111111110000110001;
		14'b00111101011010:	sigmoid = 21'b111111111110000110011;
		14'b00111101011011:	sigmoid = 21'b111111111110000110101;
		14'b00111101011100:	sigmoid = 21'b111111111110000110111;
		14'b00111101011101:	sigmoid = 21'b111111111110000111001;
		14'b00111101011110:	sigmoid = 21'b111111111110000111011;
		14'b00111101011111:	sigmoid = 21'b111111111110000111100;
		14'b00111101100000:	sigmoid = 21'b111111111110000111110;
		14'b00111101100001:	sigmoid = 21'b111111111110001000000;
		14'b00111101100010:	sigmoid = 21'b111111111110001000010;
		14'b00111101100011:	sigmoid = 21'b111111111110001000100;
		14'b00111101100100:	sigmoid = 21'b111111111110001000110;
		14'b00111101100101:	sigmoid = 21'b111111111110001001000;
		14'b00111101100110:	sigmoid = 21'b111111111110001001010;
		14'b00111101100111:	sigmoid = 21'b111111111110001001011;
		14'b00111101101000:	sigmoid = 21'b111111111110001001101;
		14'b00111101101001:	sigmoid = 21'b111111111110001001111;
		14'b00111101101010:	sigmoid = 21'b111111111110001010001;
		14'b00111101101011:	sigmoid = 21'b111111111110001010011;
		14'b00111101101100:	sigmoid = 21'b111111111110001010101;
		14'b00111101101101:	sigmoid = 21'b111111111110001010110;
		14'b00111101101110:	sigmoid = 21'b111111111110001011000;
		14'b00111101101111:	sigmoid = 21'b111111111110001011010;
		14'b00111101110000:	sigmoid = 21'b111111111110001011100;
		14'b00111101110001:	sigmoid = 21'b111111111110001011110;
		14'b00111101110010:	sigmoid = 21'b111111111110001100000;
		14'b00111101110011:	sigmoid = 21'b111111111110001100001;
		14'b00111101110100:	sigmoid = 21'b111111111110001100011;
		14'b00111101110101:	sigmoid = 21'b111111111110001100101;
		14'b00111101110110:	sigmoid = 21'b111111111110001100111;
		14'b00111101110111:	sigmoid = 21'b111111111110001101001;
		14'b00111101111000:	sigmoid = 21'b111111111110001101010;
		14'b00111101111001:	sigmoid = 21'b111111111110001101100;
		14'b00111101111010:	sigmoid = 21'b111111111110001101110;
		14'b00111101111011:	sigmoid = 21'b111111111110001110000;
		14'b00111101111100:	sigmoid = 21'b111111111110001110001;
		14'b00111101111101:	sigmoid = 21'b111111111110001110011;
		14'b00111101111110:	sigmoid = 21'b111111111110001110101;
		14'b00111101111111:	sigmoid = 21'b111111111110001110111;
		14'b00111110000000:	sigmoid = 21'b111111111110001111001;
		14'b00111110000001:	sigmoid = 21'b111111111110001111010;
		14'b00111110000010:	sigmoid = 21'b111111111110001111100;
		14'b00111110000011:	sigmoid = 21'b111111111110001111110;
		14'b00111110000100:	sigmoid = 21'b111111111110010000000;
		14'b00111110000101:	sigmoid = 21'b111111111110010000001;
		14'b00111110000110:	sigmoid = 21'b111111111110010000011;
		14'b00111110000111:	sigmoid = 21'b111111111110010000101;
		14'b00111110001000:	sigmoid = 21'b111111111110010000111;
		14'b00111110001001:	sigmoid = 21'b111111111110010001000;
		14'b00111110001010:	sigmoid = 21'b111111111110010001010;
		14'b00111110001011:	sigmoid = 21'b111111111110010001100;
		14'b00111110001100:	sigmoid = 21'b111111111110010001101;
		14'b00111110001101:	sigmoid = 21'b111111111110010001111;
		14'b00111110001110:	sigmoid = 21'b111111111110010010001;
		14'b00111110001111:	sigmoid = 21'b111111111110010010011;
		14'b00111110010000:	sigmoid = 21'b111111111110010010100;
		14'b00111110010001:	sigmoid = 21'b111111111110010010110;
		14'b00111110010010:	sigmoid = 21'b111111111110010011000;
		14'b00111110010011:	sigmoid = 21'b111111111110010011001;
		14'b00111110010100:	sigmoid = 21'b111111111110010011011;
		14'b00111110010101:	sigmoid = 21'b111111111110010011101;
		14'b00111110010110:	sigmoid = 21'b111111111110010011111;
		14'b00111110010111:	sigmoid = 21'b111111111110010100000;
		14'b00111110011000:	sigmoid = 21'b111111111110010100010;
		14'b00111110011001:	sigmoid = 21'b111111111110010100100;
		14'b00111110011010:	sigmoid = 21'b111111111110010100101;
		14'b00111110011011:	sigmoid = 21'b111111111110010100111;
		14'b00111110011100:	sigmoid = 21'b111111111110010101001;
		14'b00111110011101:	sigmoid = 21'b111111111110010101010;
		14'b00111110011110:	sigmoid = 21'b111111111110010101100;
		14'b00111110011111:	sigmoid = 21'b111111111110010101110;
		14'b00111110100000:	sigmoid = 21'b111111111110010101111;
		14'b00111110100001:	sigmoid = 21'b111111111110010110001;
		14'b00111110100010:	sigmoid = 21'b111111111110010110011;
		14'b00111110100011:	sigmoid = 21'b111111111110010110100;
		14'b00111110100100:	sigmoid = 21'b111111111110010110110;
		14'b00111110100101:	sigmoid = 21'b111111111110010110111;
		14'b00111110100110:	sigmoid = 21'b111111111110010111001;
		14'b00111110100111:	sigmoid = 21'b111111111110010111011;
		14'b00111110101000:	sigmoid = 21'b111111111110010111100;
		14'b00111110101001:	sigmoid = 21'b111111111110010111110;
		14'b00111110101010:	sigmoid = 21'b111111111110011000000;
		14'b00111110101011:	sigmoid = 21'b111111111110011000001;
		14'b00111110101100:	sigmoid = 21'b111111111110011000011;
		14'b00111110101101:	sigmoid = 21'b111111111110011000100;
		14'b00111110101110:	sigmoid = 21'b111111111110011000110;
		14'b00111110101111:	sigmoid = 21'b111111111110011001000;
		14'b00111110110000:	sigmoid = 21'b111111111110011001001;
		14'b00111110110001:	sigmoid = 21'b111111111110011001011;
		14'b00111110110010:	sigmoid = 21'b111111111110011001101;
		14'b00111110110011:	sigmoid = 21'b111111111110011001110;
		14'b00111110110100:	sigmoid = 21'b111111111110011010000;
		14'b00111110110101:	sigmoid = 21'b111111111110011010001;
		14'b00111110110110:	sigmoid = 21'b111111111110011010011;
		14'b00111110110111:	sigmoid = 21'b111111111110011010100;
		14'b00111110111000:	sigmoid = 21'b111111111110011010110;
		14'b00111110111001:	sigmoid = 21'b111111111110011011000;
		14'b00111110111010:	sigmoid = 21'b111111111110011011001;
		14'b00111110111011:	sigmoid = 21'b111111111110011011011;
		14'b00111110111100:	sigmoid = 21'b111111111110011011100;
		14'b00111110111101:	sigmoid = 21'b111111111110011011110;
		14'b00111110111110:	sigmoid = 21'b111111111110011011111;
		14'b00111110111111:	sigmoid = 21'b111111111110011100001;
		14'b00111111000000:	sigmoid = 21'b111111111110011100011;
		14'b00111111000001:	sigmoid = 21'b111111111110011100100;
		14'b00111111000010:	sigmoid = 21'b111111111110011100110;
		14'b00111111000011:	sigmoid = 21'b111111111110011100111;
		14'b00111111000100:	sigmoid = 21'b111111111110011101001;
		14'b00111111000101:	sigmoid = 21'b111111111110011101010;
		14'b00111111000110:	sigmoid = 21'b111111111110011101100;
		14'b00111111000111:	sigmoid = 21'b111111111110011101101;
		14'b00111111001000:	sigmoid = 21'b111111111110011101111;
		14'b00111111001001:	sigmoid = 21'b111111111110011110000;
		14'b00111111001010:	sigmoid = 21'b111111111110011110010;
		14'b00111111001011:	sigmoid = 21'b111111111110011110100;
		14'b00111111001100:	sigmoid = 21'b111111111110011110101;
		14'b00111111001101:	sigmoid = 21'b111111111110011110111;
		14'b00111111001110:	sigmoid = 21'b111111111110011111000;
		14'b00111111001111:	sigmoid = 21'b111111111110011111010;
		14'b00111111010000:	sigmoid = 21'b111111111110011111011;
		14'b00111111010001:	sigmoid = 21'b111111111110011111101;
		14'b00111111010010:	sigmoid = 21'b111111111110011111110;
		14'b00111111010011:	sigmoid = 21'b111111111110100000000;
		14'b00111111010100:	sigmoid = 21'b111111111110100000001;
		14'b00111111010101:	sigmoid = 21'b111111111110100000011;
		14'b00111111010110:	sigmoid = 21'b111111111110100000100;
		14'b00111111010111:	sigmoid = 21'b111111111110100000110;
		14'b00111111011000:	sigmoid = 21'b111111111110100000111;
		14'b00111111011001:	sigmoid = 21'b111111111110100001001;
		14'b00111111011010:	sigmoid = 21'b111111111110100001010;
		14'b00111111011011:	sigmoid = 21'b111111111110100001100;
		14'b00111111011100:	sigmoid = 21'b111111111110100001101;
		14'b00111111011101:	sigmoid = 21'b111111111110100001110;
		14'b00111111011110:	sigmoid = 21'b111111111110100010000;
		14'b00111111011111:	sigmoid = 21'b111111111110100010001;
		14'b00111111100000:	sigmoid = 21'b111111111110100010011;
		14'b00111111100001:	sigmoid = 21'b111111111110100010100;
		14'b00111111100010:	sigmoid = 21'b111111111110100010110;
		14'b00111111100011:	sigmoid = 21'b111111111110100010111;
		14'b00111111100100:	sigmoid = 21'b111111111110100011001;
		14'b00111111100101:	sigmoid = 21'b111111111110100011010;
		14'b00111111100110:	sigmoid = 21'b111111111110100011100;
		14'b00111111100111:	sigmoid = 21'b111111111110100011101;
		14'b00111111101000:	sigmoid = 21'b111111111110100011110;
		14'b00111111101001:	sigmoid = 21'b111111111110100100000;
		14'b00111111101010:	sigmoid = 21'b111111111110100100001;
		14'b00111111101011:	sigmoid = 21'b111111111110100100011;
		14'b00111111101100:	sigmoid = 21'b111111111110100100100;
		14'b00111111101101:	sigmoid = 21'b111111111110100100110;
		14'b00111111101110:	sigmoid = 21'b111111111110100100111;
		14'b00111111101111:	sigmoid = 21'b111111111110100101000;
		14'b00111111110000:	sigmoid = 21'b111111111110100101010;
		14'b00111111110001:	sigmoid = 21'b111111111110100101011;
		14'b00111111110010:	sigmoid = 21'b111111111110100101101;
		14'b00111111110011:	sigmoid = 21'b111111111110100101110;
		14'b00111111110100:	sigmoid = 21'b111111111110100110000;
		14'b00111111110101:	sigmoid = 21'b111111111110100110001;
		14'b00111111110110:	sigmoid = 21'b111111111110100110010;
		14'b00111111110111:	sigmoid = 21'b111111111110100110100;
		14'b00111111111000:	sigmoid = 21'b111111111110100110101;
		14'b00111111111001:	sigmoid = 21'b111111111110100110111;
		14'b00111111111010:	sigmoid = 21'b111111111110100111000;
		14'b00111111111011:	sigmoid = 21'b111111111110100111001;
		14'b00111111111100:	sigmoid = 21'b111111111110100111011;
		14'b00111111111101:	sigmoid = 21'b111111111110100111100;
		14'b00111111111110:	sigmoid = 21'b111111111110100111101;
		14'b00111111111111:	sigmoid = 21'b111111111110100111111;
		14'b01000000000000:	sigmoid = 21'b111111111110101000000;
		14'b01000000000001:	sigmoid = 21'b111111111110101000010;
		14'b01000000000010:	sigmoid = 21'b111111111110101000011;
		14'b01000000000011:	sigmoid = 21'b111111111110101000100;
		14'b01000000000100:	sigmoid = 21'b111111111110101000110;
		14'b01000000000101:	sigmoid = 21'b111111111110101000111;
		14'b01000000000110:	sigmoid = 21'b111111111110101001000;
		14'b01000000000111:	sigmoid = 21'b111111111110101001010;
		14'b01000000001000:	sigmoid = 21'b111111111110101001011;
		14'b01000000001001:	sigmoid = 21'b111111111110101001100;
		14'b01000000001010:	sigmoid = 21'b111111111110101001110;
		14'b01000000001011:	sigmoid = 21'b111111111110101001111;
		14'b01000000001100:	sigmoid = 21'b111111111110101010001;
		14'b01000000001101:	sigmoid = 21'b111111111110101010010;
		14'b01000000001110:	sigmoid = 21'b111111111110101010011;
		14'b01000000001111:	sigmoid = 21'b111111111110101010101;
		14'b01000000010000:	sigmoid = 21'b111111111110101010110;
		14'b01000000010001:	sigmoid = 21'b111111111110101010111;
		14'b01000000010010:	sigmoid = 21'b111111111110101011001;
		14'b01000000010011:	sigmoid = 21'b111111111110101011010;
		14'b01000000010100:	sigmoid = 21'b111111111110101011011;
		14'b01000000010101:	sigmoid = 21'b111111111110101011100;
		14'b01000000010110:	sigmoid = 21'b111111111110101011110;
		14'b01000000010111:	sigmoid = 21'b111111111110101011111;
		14'b01000000011000:	sigmoid = 21'b111111111110101100000;
		14'b01000000011001:	sigmoid = 21'b111111111110101100010;
		14'b01000000011010:	sigmoid = 21'b111111111110101100011;
		14'b01000000011011:	sigmoid = 21'b111111111110101100100;
		14'b01000000011100:	sigmoid = 21'b111111111110101100110;
		14'b01000000011101:	sigmoid = 21'b111111111110101100111;
		14'b01000000011110:	sigmoid = 21'b111111111110101101000;
		14'b01000000011111:	sigmoid = 21'b111111111110101101010;
		14'b01000000100000:	sigmoid = 21'b111111111110101101011;
		14'b01000000100001:	sigmoid = 21'b111111111110101101100;
		14'b01000000100010:	sigmoid = 21'b111111111110101101101;
		14'b01000000100011:	sigmoid = 21'b111111111110101101111;
		14'b01000000100100:	sigmoid = 21'b111111111110101110000;
		14'b01000000100101:	sigmoid = 21'b111111111110101110001;
		14'b01000000100110:	sigmoid = 21'b111111111110101110011;
		14'b01000000100111:	sigmoid = 21'b111111111110101110100;
		14'b01000000101000:	sigmoid = 21'b111111111110101110101;
		14'b01000000101001:	sigmoid = 21'b111111111110101110110;
		14'b01000000101010:	sigmoid = 21'b111111111110101111000;
		14'b01000000101011:	sigmoid = 21'b111111111110101111001;
		14'b01000000101100:	sigmoid = 21'b111111111110101111010;
		14'b01000000101101:	sigmoid = 21'b111111111110101111011;
		14'b01000000101110:	sigmoid = 21'b111111111110101111101;
		14'b01000000101111:	sigmoid = 21'b111111111110101111110;
		14'b01000000110000:	sigmoid = 21'b111111111110101111111;
		14'b01000000110001:	sigmoid = 21'b111111111110110000000;
		14'b01000000110010:	sigmoid = 21'b111111111110110000010;
		14'b01000000110011:	sigmoid = 21'b111111111110110000011;
		14'b01000000110100:	sigmoid = 21'b111111111110110000100;
		14'b01000000110101:	sigmoid = 21'b111111111110110000101;
		14'b01000000110110:	sigmoid = 21'b111111111110110000111;
		14'b01000000110111:	sigmoid = 21'b111111111110110001000;
		14'b01000000111000:	sigmoid = 21'b111111111110110001001;
		14'b01000000111001:	sigmoid = 21'b111111111110110001010;
		14'b01000000111010:	sigmoid = 21'b111111111110110001100;
		14'b01000000111011:	sigmoid = 21'b111111111110110001101;
		14'b01000000111100:	sigmoid = 21'b111111111110110001110;
		14'b01000000111101:	sigmoid = 21'b111111111110110001111;
		14'b01000000111110:	sigmoid = 21'b111111111110110010000;
		14'b01000000111111:	sigmoid = 21'b111111111110110010010;
		14'b01000001000000:	sigmoid = 21'b111111111110110010011;
		14'b01000001000001:	sigmoid = 21'b111111111110110010100;
		14'b01000001000010:	sigmoid = 21'b111111111110110010101;
		14'b01000001000011:	sigmoid = 21'b111111111110110010110;
		14'b01000001000100:	sigmoid = 21'b111111111110110011000;
		14'b01000001000101:	sigmoid = 21'b111111111110110011001;
		14'b01000001000110:	sigmoid = 21'b111111111110110011010;
		14'b01000001000111:	sigmoid = 21'b111111111110110011011;
		14'b01000001001000:	sigmoid = 21'b111111111110110011100;
		14'b01000001001001:	sigmoid = 21'b111111111110110011110;
		14'b01000001001010:	sigmoid = 21'b111111111110110011111;
		14'b01000001001011:	sigmoid = 21'b111111111110110100000;
		14'b01000001001100:	sigmoid = 21'b111111111110110100001;
		14'b01000001001101:	sigmoid = 21'b111111111110110100010;
		14'b01000001001110:	sigmoid = 21'b111111111110110100100;
		14'b01000001001111:	sigmoid = 21'b111111111110110100101;
		14'b01000001010000:	sigmoid = 21'b111111111110110100110;
		14'b01000001010001:	sigmoid = 21'b111111111110110100111;
		14'b01000001010010:	sigmoid = 21'b111111111110110101000;
		14'b01000001010011:	sigmoid = 21'b111111111110110101001;
		14'b01000001010100:	sigmoid = 21'b111111111110110101011;
		14'b01000001010101:	sigmoid = 21'b111111111110110101100;
		14'b01000001010110:	sigmoid = 21'b111111111110110101101;
		14'b01000001010111:	sigmoid = 21'b111111111110110101110;
		14'b01000001011000:	sigmoid = 21'b111111111110110101111;
		14'b01000001011001:	sigmoid = 21'b111111111110110110000;
		14'b01000001011010:	sigmoid = 21'b111111111110110110010;
		14'b01000001011011:	sigmoid = 21'b111111111110110110011;
		14'b01000001011100:	sigmoid = 21'b111111111110110110100;
		14'b01000001011101:	sigmoid = 21'b111111111110110110101;
		14'b01000001011110:	sigmoid = 21'b111111111110110110110;
		14'b01000001011111:	sigmoid = 21'b111111111110110110111;
		14'b01000001100000:	sigmoid = 21'b111111111110110111000;
		14'b01000001100001:	sigmoid = 21'b111111111110110111010;
		14'b01000001100010:	sigmoid = 21'b111111111110110111011;
		14'b01000001100011:	sigmoid = 21'b111111111110110111100;
		14'b01000001100100:	sigmoid = 21'b111111111110110111101;
		14'b01000001100101:	sigmoid = 21'b111111111110110111110;
		14'b01000001100110:	sigmoid = 21'b111111111110110111111;
		14'b01000001100111:	sigmoid = 21'b111111111110111000000;
		14'b01000001101000:	sigmoid = 21'b111111111110111000001;
		14'b01000001101001:	sigmoid = 21'b111111111110111000011;
		14'b01000001101010:	sigmoid = 21'b111111111110111000100;
		14'b01000001101011:	sigmoid = 21'b111111111110111000101;
		14'b01000001101100:	sigmoid = 21'b111111111110111000110;
		14'b01000001101101:	sigmoid = 21'b111111111110111000111;
		14'b01000001101110:	sigmoid = 21'b111111111110111001000;
		14'b01000001101111:	sigmoid = 21'b111111111110111001001;
		14'b01000001110000:	sigmoid = 21'b111111111110111001010;
		14'b01000001110001:	sigmoid = 21'b111111111110111001011;
		14'b01000001110010:	sigmoid = 21'b111111111110111001101;
		14'b01000001110011:	sigmoid = 21'b111111111110111001110;
		14'b01000001110100:	sigmoid = 21'b111111111110111001111;
		14'b01000001110101:	sigmoid = 21'b111111111110111010000;
		14'b01000001110110:	sigmoid = 21'b111111111110111010001;
		14'b01000001110111:	sigmoid = 21'b111111111110111010010;
		14'b01000001111000:	sigmoid = 21'b111111111110111010011;
		14'b01000001111001:	sigmoid = 21'b111111111110111010100;
		14'b01000001111010:	sigmoid = 21'b111111111110111010101;
		14'b01000001111011:	sigmoid = 21'b111111111110111010110;
		14'b01000001111100:	sigmoid = 21'b111111111110111010111;
		14'b01000001111101:	sigmoid = 21'b111111111110111011001;
		14'b01000001111110:	sigmoid = 21'b111111111110111011010;
		14'b01000001111111:	sigmoid = 21'b111111111110111011011;
		14'b01000010000000:	sigmoid = 21'b111111111110111011100;
		14'b01000010000001:	sigmoid = 21'b111111111110111011101;
		14'b01000010000010:	sigmoid = 21'b111111111110111011110;
		14'b01000010000011:	sigmoid = 21'b111111111110111011111;
		14'b01000010000100:	sigmoid = 21'b111111111110111100000;
		14'b01000010000101:	sigmoid = 21'b111111111110111100001;
		14'b01000010000110:	sigmoid = 21'b111111111110111100010;
		14'b01000010000111:	sigmoid = 21'b111111111110111100011;
		14'b01000010001000:	sigmoid = 21'b111111111110111100100;
		14'b01000010001001:	sigmoid = 21'b111111111110111100101;
		14'b01000010001010:	sigmoid = 21'b111111111110111100110;
		14'b01000010001011:	sigmoid = 21'b111111111110111100111;
		14'b01000010001100:	sigmoid = 21'b111111111110111101000;
		14'b01000010001101:	sigmoid = 21'b111111111110111101001;
		14'b01000010001110:	sigmoid = 21'b111111111110111101011;
		14'b01000010001111:	sigmoid = 21'b111111111110111101100;
		14'b01000010010000:	sigmoid = 21'b111111111110111101101;
		14'b01000010010001:	sigmoid = 21'b111111111110111101110;
		14'b01000010010010:	sigmoid = 21'b111111111110111101111;
		14'b01000010010011:	sigmoid = 21'b111111111110111110000;
		14'b01000010010100:	sigmoid = 21'b111111111110111110001;
		14'b01000010010101:	sigmoid = 21'b111111111110111110010;
		14'b01000010010110:	sigmoid = 21'b111111111110111110011;
		14'b01000010010111:	sigmoid = 21'b111111111110111110100;
		14'b01000010011000:	sigmoid = 21'b111111111110111110101;
		14'b01000010011001:	sigmoid = 21'b111111111110111110110;
		14'b01000010011010:	sigmoid = 21'b111111111110111110111;
		14'b01000010011011:	sigmoid = 21'b111111111110111111000;
		14'b01000010011100:	sigmoid = 21'b111111111110111111001;
		14'b01000010011101:	sigmoid = 21'b111111111110111111010;
		14'b01000010011110:	sigmoid = 21'b111111111110111111011;
		14'b01000010011111:	sigmoid = 21'b111111111110111111100;
		14'b01000010100000:	sigmoid = 21'b111111111110111111101;
		14'b01000010100001:	sigmoid = 21'b111111111110111111110;
		14'b01000010100010:	sigmoid = 21'b111111111110111111111;
		14'b01000010100011:	sigmoid = 21'b111111111111000000000;
		14'b01000010100100:	sigmoid = 21'b111111111111000000001;
		14'b01000010100101:	sigmoid = 21'b111111111111000000010;
		14'b01000010100110:	sigmoid = 21'b111111111111000000011;
		14'b01000010100111:	sigmoid = 21'b111111111111000000100;
		14'b01000010101000:	sigmoid = 21'b111111111111000000101;
		14'b01000010101001:	sigmoid = 21'b111111111111000000110;
		14'b01000010101010:	sigmoid = 21'b111111111111000000111;
		14'b01000010101011:	sigmoid = 21'b111111111111000001000;
		14'b01000010101100:	sigmoid = 21'b111111111111000001001;
		14'b01000010101101:	sigmoid = 21'b111111111111000001010;
		14'b01000010101110:	sigmoid = 21'b111111111111000001011;
		14'b01000010101111:	sigmoid = 21'b111111111111000001100;
		14'b01000010110000:	sigmoid = 21'b111111111111000001101;
		14'b01000010110001:	sigmoid = 21'b111111111111000001110;
		14'b01000010110010:	sigmoid = 21'b111111111111000001111;
		14'b01000010110011:	sigmoid = 21'b111111111111000010000;
		14'b01000010110100:	sigmoid = 21'b111111111111000010001;
		14'b01000010110101:	sigmoid = 21'b111111111111000010010;
		14'b01000010110110:	sigmoid = 21'b111111111111000010011;
		14'b01000010110111:	sigmoid = 21'b111111111111000010100;
		14'b01000010111000:	sigmoid = 21'b111111111111000010100;
		14'b01000010111001:	sigmoid = 21'b111111111111000010101;
		14'b01000010111010:	sigmoid = 21'b111111111111000010110;
		14'b01000010111011:	sigmoid = 21'b111111111111000010111;
		14'b01000010111100:	sigmoid = 21'b111111111111000011000;
		14'b01000010111101:	sigmoid = 21'b111111111111000011001;
		14'b01000010111110:	sigmoid = 21'b111111111111000011010;
		14'b01000010111111:	sigmoid = 21'b111111111111000011011;
		14'b01000011000000:	sigmoid = 21'b111111111111000011100;
		14'b01000011000001:	sigmoid = 21'b111111111111000011101;
		14'b01000011000010:	sigmoid = 21'b111111111111000011110;
		14'b01000011000011:	sigmoid = 21'b111111111111000011111;
		14'b01000011000100:	sigmoid = 21'b111111111111000100000;
		14'b01000011000101:	sigmoid = 21'b111111111111000100001;
		14'b01000011000110:	sigmoid = 21'b111111111111000100010;
		14'b01000011000111:	sigmoid = 21'b111111111111000100011;
		14'b01000011001000:	sigmoid = 21'b111111111111000100100;
		14'b01000011001001:	sigmoid = 21'b111111111111000100101;
		14'b01000011001010:	sigmoid = 21'b111111111111000100101;
		14'b01000011001011:	sigmoid = 21'b111111111111000100110;
		14'b01000011001100:	sigmoid = 21'b111111111111000100111;
		14'b01000011001101:	sigmoid = 21'b111111111111000101000;
		14'b01000011001110:	sigmoid = 21'b111111111111000101001;
		14'b01000011001111:	sigmoid = 21'b111111111111000101010;
		14'b01000011010000:	sigmoid = 21'b111111111111000101011;
		14'b01000011010001:	sigmoid = 21'b111111111111000101100;
		14'b01000011010010:	sigmoid = 21'b111111111111000101101;
		14'b01000011010011:	sigmoid = 21'b111111111111000101110;
		14'b01000011010100:	sigmoid = 21'b111111111111000101111;
		14'b01000011010101:	sigmoid = 21'b111111111111000110000;
		14'b01000011010110:	sigmoid = 21'b111111111111000110000;
		14'b01000011010111:	sigmoid = 21'b111111111111000110001;
		14'b01000011011000:	sigmoid = 21'b111111111111000110010;
		14'b01000011011001:	sigmoid = 21'b111111111111000110011;
		14'b01000011011010:	sigmoid = 21'b111111111111000110100;
		14'b01000011011011:	sigmoid = 21'b111111111111000110101;
		14'b01000011011100:	sigmoid = 21'b111111111111000110110;
		14'b01000011011101:	sigmoid = 21'b111111111111000110111;
		14'b01000011011110:	sigmoid = 21'b111111111111000111000;
		14'b01000011011111:	sigmoid = 21'b111111111111000111000;
		14'b01000011100000:	sigmoid = 21'b111111111111000111001;
		14'b01000011100001:	sigmoid = 21'b111111111111000111010;
		14'b01000011100010:	sigmoid = 21'b111111111111000111011;
		14'b01000011100011:	sigmoid = 21'b111111111111000111100;
		14'b01000011100100:	sigmoid = 21'b111111111111000111101;
		14'b01000011100101:	sigmoid = 21'b111111111111000111110;
		14'b01000011100110:	sigmoid = 21'b111111111111000111111;
		14'b01000011100111:	sigmoid = 21'b111111111111001000000;
		14'b01000011101000:	sigmoid = 21'b111111111111001000000;
		14'b01000011101001:	sigmoid = 21'b111111111111001000001;
		14'b01000011101010:	sigmoid = 21'b111111111111001000010;
		14'b01000011101011:	sigmoid = 21'b111111111111001000011;
		14'b01000011101100:	sigmoid = 21'b111111111111001000100;
		14'b01000011101101:	sigmoid = 21'b111111111111001000101;
		14'b01000011101110:	sigmoid = 21'b111111111111001000110;
		14'b01000011101111:	sigmoid = 21'b111111111111001000110;
		14'b01000011110000:	sigmoid = 21'b111111111111001000111;
		14'b01000011110001:	sigmoid = 21'b111111111111001001000;
		14'b01000011110010:	sigmoid = 21'b111111111111001001001;
		14'b01000011110011:	sigmoid = 21'b111111111111001001010;
		14'b01000011110100:	sigmoid = 21'b111111111111001001011;
		14'b01000011110101:	sigmoid = 21'b111111111111001001100;
		14'b01000011110110:	sigmoid = 21'b111111111111001001100;
		14'b01000011110111:	sigmoid = 21'b111111111111001001101;
		14'b01000011111000:	sigmoid = 21'b111111111111001001110;
		14'b01000011111001:	sigmoid = 21'b111111111111001001111;
		14'b01000011111010:	sigmoid = 21'b111111111111001010000;
		14'b01000011111011:	sigmoid = 21'b111111111111001010001;
		14'b01000011111100:	sigmoid = 21'b111111111111001010010;
		14'b01000011111101:	sigmoid = 21'b111111111111001010010;
		14'b01000011111110:	sigmoid = 21'b111111111111001010011;
		14'b01000011111111:	sigmoid = 21'b111111111111001010100;
		14'b01000100000000:	sigmoid = 21'b111111111111001010101;
		14'b01000100000001:	sigmoid = 21'b111111111111001010110;
		14'b01000100000010:	sigmoid = 21'b111111111111001010111;
		14'b01000100000011:	sigmoid = 21'b111111111111001010111;
		14'b01000100000100:	sigmoid = 21'b111111111111001011000;
		14'b01000100000101:	sigmoid = 21'b111111111111001011001;
		14'b01000100000110:	sigmoid = 21'b111111111111001011010;
		14'b01000100000111:	sigmoid = 21'b111111111111001011011;
		14'b01000100001000:	sigmoid = 21'b111111111111001011011;
		14'b01000100001001:	sigmoid = 21'b111111111111001011100;
		14'b01000100001010:	sigmoid = 21'b111111111111001011101;
		14'b01000100001011:	sigmoid = 21'b111111111111001011110;
		14'b01000100001100:	sigmoid = 21'b111111111111001011111;
		14'b01000100001101:	sigmoid = 21'b111111111111001100000;
		14'b01000100001110:	sigmoid = 21'b111111111111001100000;
		14'b01000100001111:	sigmoid = 21'b111111111111001100001;
		14'b01000100010000:	sigmoid = 21'b111111111111001100010;
		14'b01000100010001:	sigmoid = 21'b111111111111001100011;
		14'b01000100010010:	sigmoid = 21'b111111111111001100100;
		14'b01000100010011:	sigmoid = 21'b111111111111001100100;
		14'b01000100010100:	sigmoid = 21'b111111111111001100101;
		14'b01000100010101:	sigmoid = 21'b111111111111001100110;
		14'b01000100010110:	sigmoid = 21'b111111111111001100111;
		14'b01000100010111:	sigmoid = 21'b111111111111001101000;
		14'b01000100011000:	sigmoid = 21'b111111111111001101000;
		14'b01000100011001:	sigmoid = 21'b111111111111001101001;
		14'b01000100011010:	sigmoid = 21'b111111111111001101010;
		14'b01000100011011:	sigmoid = 21'b111111111111001101011;
		14'b01000100011100:	sigmoid = 21'b111111111111001101100;
		14'b01000100011101:	sigmoid = 21'b111111111111001101100;
		14'b01000100011110:	sigmoid = 21'b111111111111001101101;
		14'b01000100011111:	sigmoid = 21'b111111111111001101110;
		14'b01000100100000:	sigmoid = 21'b111111111111001101111;
		14'b01000100100001:	sigmoid = 21'b111111111111001110000;
		14'b01000100100010:	sigmoid = 21'b111111111111001110000;
		14'b01000100100011:	sigmoid = 21'b111111111111001110001;
		14'b01000100100100:	sigmoid = 21'b111111111111001110010;
		14'b01000100100101:	sigmoid = 21'b111111111111001110011;
		14'b01000100100110:	sigmoid = 21'b111111111111001110011;
		14'b01000100100111:	sigmoid = 21'b111111111111001110100;
		14'b01000100101000:	sigmoid = 21'b111111111111001110101;
		14'b01000100101001:	sigmoid = 21'b111111111111001110110;
		14'b01000100101010:	sigmoid = 21'b111111111111001110110;
		14'b01000100101011:	sigmoid = 21'b111111111111001110111;
		14'b01000100101100:	sigmoid = 21'b111111111111001111000;
		14'b01000100101101:	sigmoid = 21'b111111111111001111001;
		14'b01000100101110:	sigmoid = 21'b111111111111001111010;
		14'b01000100101111:	sigmoid = 21'b111111111111001111010;
		14'b01000100110000:	sigmoid = 21'b111111111111001111011;
		14'b01000100110001:	sigmoid = 21'b111111111111001111100;
		14'b01000100110010:	sigmoid = 21'b111111111111001111101;
		14'b01000100110011:	sigmoid = 21'b111111111111001111101;
		14'b01000100110100:	sigmoid = 21'b111111111111001111110;
		14'b01000100110101:	sigmoid = 21'b111111111111001111111;
		14'b01000100110110:	sigmoid = 21'b111111111111010000000;
		14'b01000100110111:	sigmoid = 21'b111111111111010000000;
		14'b01000100111000:	sigmoid = 21'b111111111111010000001;
		14'b01000100111001:	sigmoid = 21'b111111111111010000010;
		14'b01000100111010:	sigmoid = 21'b111111111111010000011;
		14'b01000100111011:	sigmoid = 21'b111111111111010000011;
		14'b01000100111100:	sigmoid = 21'b111111111111010000100;
		14'b01000100111101:	sigmoid = 21'b111111111111010000101;
		14'b01000100111110:	sigmoid = 21'b111111111111010000110;
		14'b01000100111111:	sigmoid = 21'b111111111111010000110;
		14'b01000101000000:	sigmoid = 21'b111111111111010000111;
		14'b01000101000001:	sigmoid = 21'b111111111111010001000;
		14'b01000101000010:	sigmoid = 21'b111111111111010001000;
		14'b01000101000011:	sigmoid = 21'b111111111111010001001;
		14'b01000101000100:	sigmoid = 21'b111111111111010001010;
		14'b01000101000101:	sigmoid = 21'b111111111111010001011;
		14'b01000101000110:	sigmoid = 21'b111111111111010001011;
		14'b01000101000111:	sigmoid = 21'b111111111111010001100;
		14'b01000101001000:	sigmoid = 21'b111111111111010001101;
		14'b01000101001001:	sigmoid = 21'b111111111111010001110;
		14'b01000101001010:	sigmoid = 21'b111111111111010001110;
		14'b01000101001011:	sigmoid = 21'b111111111111010001111;
		14'b01000101001100:	sigmoid = 21'b111111111111010010000;
		14'b01000101001101:	sigmoid = 21'b111111111111010010000;
		14'b01000101001110:	sigmoid = 21'b111111111111010010001;
		14'b01000101001111:	sigmoid = 21'b111111111111010010010;
		14'b01000101010000:	sigmoid = 21'b111111111111010010011;
		14'b01000101010001:	sigmoid = 21'b111111111111010010011;
		14'b01000101010010:	sigmoid = 21'b111111111111010010100;
		14'b01000101010011:	sigmoid = 21'b111111111111010010101;
		14'b01000101010100:	sigmoid = 21'b111111111111010010101;
		14'b01000101010101:	sigmoid = 21'b111111111111010010110;
		14'b01000101010110:	sigmoid = 21'b111111111111010010111;
		14'b01000101010111:	sigmoid = 21'b111111111111010011000;
		14'b01000101011000:	sigmoid = 21'b111111111111010011000;
		14'b01000101011001:	sigmoid = 21'b111111111111010011001;
		14'b01000101011010:	sigmoid = 21'b111111111111010011010;
		14'b01000101011011:	sigmoid = 21'b111111111111010011010;
		14'b01000101011100:	sigmoid = 21'b111111111111010011011;
		14'b01000101011101:	sigmoid = 21'b111111111111010011100;
		14'b01000101011110:	sigmoid = 21'b111111111111010011100;
		14'b01000101011111:	sigmoid = 21'b111111111111010011101;
		14'b01000101100000:	sigmoid = 21'b111111111111010011110;
		14'b01000101100001:	sigmoid = 21'b111111111111010011110;
		14'b01000101100010:	sigmoid = 21'b111111111111010011111;
		14'b01000101100011:	sigmoid = 21'b111111111111010100000;
		14'b01000101100100:	sigmoid = 21'b111111111111010100001;
		14'b01000101100101:	sigmoid = 21'b111111111111010100001;
		14'b01000101100110:	sigmoid = 21'b111111111111010100010;
		14'b01000101100111:	sigmoid = 21'b111111111111010100011;
		14'b01000101101000:	sigmoid = 21'b111111111111010100011;
		14'b01000101101001:	sigmoid = 21'b111111111111010100100;
		14'b01000101101010:	sigmoid = 21'b111111111111010100101;
		14'b01000101101011:	sigmoid = 21'b111111111111010100101;
		14'b01000101101100:	sigmoid = 21'b111111111111010100110;
		14'b01000101101101:	sigmoid = 21'b111111111111010100111;
		14'b01000101101110:	sigmoid = 21'b111111111111010100111;
		14'b01000101101111:	sigmoid = 21'b111111111111010101000;
		14'b01000101110000:	sigmoid = 21'b111111111111010101001;
		14'b01000101110001:	sigmoid = 21'b111111111111010101001;
		14'b01000101110010:	sigmoid = 21'b111111111111010101010;
		14'b01000101110011:	sigmoid = 21'b111111111111010101011;
		14'b01000101110100:	sigmoid = 21'b111111111111010101011;
		14'b01000101110101:	sigmoid = 21'b111111111111010101100;
		14'b01000101110110:	sigmoid = 21'b111111111111010101101;
		14'b01000101110111:	sigmoid = 21'b111111111111010101101;
		14'b01000101111000:	sigmoid = 21'b111111111111010101110;
		14'b01000101111001:	sigmoid = 21'b111111111111010101111;
		14'b01000101111010:	sigmoid = 21'b111111111111010101111;
		14'b01000101111011:	sigmoid = 21'b111111111111010110000;
		14'b01000101111100:	sigmoid = 21'b111111111111010110001;
		14'b01000101111101:	sigmoid = 21'b111111111111010110001;
		14'b01000101111110:	sigmoid = 21'b111111111111010110010;
		14'b01000101111111:	sigmoid = 21'b111111111111010110011;
		14'b01000110000000:	sigmoid = 21'b111111111111010110011;
		14'b01000110000001:	sigmoid = 21'b111111111111010110100;
		14'b01000110000010:	sigmoid = 21'b111111111111010110101;
		14'b01000110000011:	sigmoid = 21'b111111111111010110101;
		14'b01000110000100:	sigmoid = 21'b111111111111010110110;
		14'b01000110000101:	sigmoid = 21'b111111111111010110110;
		14'b01000110000110:	sigmoid = 21'b111111111111010110111;
		14'b01000110000111:	sigmoid = 21'b111111111111010111000;
		14'b01000110001000:	sigmoid = 21'b111111111111010111000;
		14'b01000110001001:	sigmoid = 21'b111111111111010111001;
		14'b01000110001010:	sigmoid = 21'b111111111111010111010;
		14'b01000110001011:	sigmoid = 21'b111111111111010111010;
		14'b01000110001100:	sigmoid = 21'b111111111111010111011;
		14'b01000110001101:	sigmoid = 21'b111111111111010111100;
		14'b01000110001110:	sigmoid = 21'b111111111111010111100;
		14'b01000110001111:	sigmoid = 21'b111111111111010111101;
		14'b01000110010000:	sigmoid = 21'b111111111111010111101;
		14'b01000110010001:	sigmoid = 21'b111111111111010111110;
		14'b01000110010010:	sigmoid = 21'b111111111111010111111;
		14'b01000110010011:	sigmoid = 21'b111111111111010111111;
		14'b01000110010100:	sigmoid = 21'b111111111111011000000;
		14'b01000110010101:	sigmoid = 21'b111111111111011000001;
		14'b01000110010110:	sigmoid = 21'b111111111111011000001;
		14'b01000110010111:	sigmoid = 21'b111111111111011000010;
		14'b01000110011000:	sigmoid = 21'b111111111111011000010;
		14'b01000110011001:	sigmoid = 21'b111111111111011000011;
		14'b01000110011010:	sigmoid = 21'b111111111111011000100;
		14'b01000110011011:	sigmoid = 21'b111111111111011000100;
		14'b01000110011100:	sigmoid = 21'b111111111111011000101;
		14'b01000110011101:	sigmoid = 21'b111111111111011000110;
		14'b01000110011110:	sigmoid = 21'b111111111111011000110;
		14'b01000110011111:	sigmoid = 21'b111111111111011000111;
		14'b01000110100000:	sigmoid = 21'b111111111111011000111;
		14'b01000110100001:	sigmoid = 21'b111111111111011001000;
		14'b01000110100010:	sigmoid = 21'b111111111111011001001;
		14'b01000110100011:	sigmoid = 21'b111111111111011001001;
		14'b01000110100100:	sigmoid = 21'b111111111111011001010;
		14'b01000110100101:	sigmoid = 21'b111111111111011001010;
		14'b01000110100110:	sigmoid = 21'b111111111111011001011;
		14'b01000110100111:	sigmoid = 21'b111111111111011001100;
		14'b01000110101000:	sigmoid = 21'b111111111111011001100;
		14'b01000110101001:	sigmoid = 21'b111111111111011001101;
		14'b01000110101010:	sigmoid = 21'b111111111111011001101;
		14'b01000110101011:	sigmoid = 21'b111111111111011001110;
		14'b01000110101100:	sigmoid = 21'b111111111111011001111;
		14'b01000110101101:	sigmoid = 21'b111111111111011001111;
		14'b01000110101110:	sigmoid = 21'b111111111111011010000;
		14'b01000110101111:	sigmoid = 21'b111111111111011010000;
		14'b01000110110000:	sigmoid = 21'b111111111111011010001;
		14'b01000110110001:	sigmoid = 21'b111111111111011010010;
		14'b01000110110010:	sigmoid = 21'b111111111111011010010;
		14'b01000110110011:	sigmoid = 21'b111111111111011010011;
		14'b01000110110100:	sigmoid = 21'b111111111111011010011;
		14'b01000110110101:	sigmoid = 21'b111111111111011010100;
		14'b01000110110110:	sigmoid = 21'b111111111111011010100;
		14'b01000110110111:	sigmoid = 21'b111111111111011010101;
		14'b01000110111000:	sigmoid = 21'b111111111111011010110;
		14'b01000110111001:	sigmoid = 21'b111111111111011010110;
		14'b01000110111010:	sigmoid = 21'b111111111111011010111;
		14'b01000110111011:	sigmoid = 21'b111111111111011010111;
		14'b01000110111100:	sigmoid = 21'b111111111111011011000;
		14'b01000110111101:	sigmoid = 21'b111111111111011011001;
		14'b01000110111110:	sigmoid = 21'b111111111111011011001;
		14'b01000110111111:	sigmoid = 21'b111111111111011011010;
		14'b01000111000000:	sigmoid = 21'b111111111111011011010;
		14'b01000111000001:	sigmoid = 21'b111111111111011011011;
		14'b01000111000010:	sigmoid = 21'b111111111111011011011;
		14'b01000111000011:	sigmoid = 21'b111111111111011011100;
		14'b01000111000100:	sigmoid = 21'b111111111111011011101;
		14'b01000111000101:	sigmoid = 21'b111111111111011011101;
		14'b01000111000110:	sigmoid = 21'b111111111111011011110;
		14'b01000111000111:	sigmoid = 21'b111111111111011011110;
		14'b01000111001000:	sigmoid = 21'b111111111111011011111;
		14'b01000111001001:	sigmoid = 21'b111111111111011011111;
		14'b01000111001010:	sigmoid = 21'b111111111111011100000;
		14'b01000111001011:	sigmoid = 21'b111111111111011100001;
		14'b01000111001100:	sigmoid = 21'b111111111111011100001;
		14'b01000111001101:	sigmoid = 21'b111111111111011100010;
		14'b01000111001110:	sigmoid = 21'b111111111111011100010;
		14'b01000111001111:	sigmoid = 21'b111111111111011100011;
		14'b01000111010000:	sigmoid = 21'b111111111111011100011;
		14'b01000111010001:	sigmoid = 21'b111111111111011100100;
		14'b01000111010010:	sigmoid = 21'b111111111111011100100;
		14'b01000111010011:	sigmoid = 21'b111111111111011100101;
		14'b01000111010100:	sigmoid = 21'b111111111111011100110;
		14'b01000111010101:	sigmoid = 21'b111111111111011100110;
		14'b01000111010110:	sigmoid = 21'b111111111111011100111;
		14'b01000111010111:	sigmoid = 21'b111111111111011100111;
		14'b01000111011000:	sigmoid = 21'b111111111111011101000;
		14'b01000111011001:	sigmoid = 21'b111111111111011101000;
		14'b01000111011010:	sigmoid = 21'b111111111111011101001;
		14'b01000111011011:	sigmoid = 21'b111111111111011101001;
		14'b01000111011100:	sigmoid = 21'b111111111111011101010;
		14'b01000111011101:	sigmoid = 21'b111111111111011101010;
		14'b01000111011110:	sigmoid = 21'b111111111111011101011;
		14'b01000111011111:	sigmoid = 21'b111111111111011101011;
		14'b01000111100000:	sigmoid = 21'b111111111111011101100;
		14'b01000111100001:	sigmoid = 21'b111111111111011101101;
		14'b01000111100010:	sigmoid = 21'b111111111111011101101;
		14'b01000111100011:	sigmoid = 21'b111111111111011101110;
		14'b01000111100100:	sigmoid = 21'b111111111111011101110;
		14'b01000111100101:	sigmoid = 21'b111111111111011101111;
		14'b01000111100110:	sigmoid = 21'b111111111111011101111;
		14'b01000111100111:	sigmoid = 21'b111111111111011110000;
		14'b01000111101000:	sigmoid = 21'b111111111111011110000;
		14'b01000111101001:	sigmoid = 21'b111111111111011110001;
		14'b01000111101010:	sigmoid = 21'b111111111111011110001;
		14'b01000111101011:	sigmoid = 21'b111111111111011110010;
		14'b01000111101100:	sigmoid = 21'b111111111111011110010;
		14'b01000111101101:	sigmoid = 21'b111111111111011110011;
		14'b01000111101110:	sigmoid = 21'b111111111111011110011;
		14'b01000111101111:	sigmoid = 21'b111111111111011110100;
		14'b01000111110000:	sigmoid = 21'b111111111111011110101;
		14'b01000111110001:	sigmoid = 21'b111111111111011110101;
		14'b01000111110010:	sigmoid = 21'b111111111111011110110;
		14'b01000111110011:	sigmoid = 21'b111111111111011110110;
		14'b01000111110100:	sigmoid = 21'b111111111111011110111;
		14'b01000111110101:	sigmoid = 21'b111111111111011110111;
		14'b01000111110110:	sigmoid = 21'b111111111111011111000;
		14'b01000111110111:	sigmoid = 21'b111111111111011111000;
		14'b01000111111000:	sigmoid = 21'b111111111111011111001;
		14'b01000111111001:	sigmoid = 21'b111111111111011111001;
		14'b01000111111010:	sigmoid = 21'b111111111111011111010;
		14'b01000111111011:	sigmoid = 21'b111111111111011111010;
		14'b01000111111100:	sigmoid = 21'b111111111111011111011;
		14'b01000111111101:	sigmoid = 21'b111111111111011111011;
		14'b01000111111110:	sigmoid = 21'b111111111111011111100;
		14'b01000111111111:	sigmoid = 21'b111111111111011111100;
		14'b01001000000000:	sigmoid = 21'b111111111111011111101;
		14'b01001000000001:	sigmoid = 21'b111111111111011111101;
		14'b01001000000010:	sigmoid = 21'b111111111111011111110;
		14'b01001000000011:	sigmoid = 21'b111111111111011111110;
		14'b01001000000100:	sigmoid = 21'b111111111111011111111;
		14'b01001000000101:	sigmoid = 21'b111111111111011111111;
		14'b01001000000110:	sigmoid = 21'b111111111111100000000;
		14'b01001000000111:	sigmoid = 21'b111111111111100000000;
		14'b01001000001000:	sigmoid = 21'b111111111111100000001;
		14'b01001000001001:	sigmoid = 21'b111111111111100000001;
		14'b01001000001010:	sigmoid = 21'b111111111111100000010;
		14'b01001000001011:	sigmoid = 21'b111111111111100000010;
		14'b01001000001100:	sigmoid = 21'b111111111111100000011;
		14'b01001000001101:	sigmoid = 21'b111111111111100000011;
		14'b01001000001110:	sigmoid = 21'b111111111111100000100;
		14'b01001000001111:	sigmoid = 21'b111111111111100000100;
		14'b01001000010000:	sigmoid = 21'b111111111111100000101;
		14'b01001000010001:	sigmoid = 21'b111111111111100000101;
		14'b01001000010010:	sigmoid = 21'b111111111111100000110;
		14'b01001000010011:	sigmoid = 21'b111111111111100000110;
		14'b01001000010100:	sigmoid = 21'b111111111111100000111;
		14'b01001000010101:	sigmoid = 21'b111111111111100000111;
		14'b01001000010110:	sigmoid = 21'b111111111111100001000;
		14'b01001000010111:	sigmoid = 21'b111111111111100001000;
		14'b01001000011000:	sigmoid = 21'b111111111111100001001;
		14'b01001000011001:	sigmoid = 21'b111111111111100001001;
		14'b01001000011010:	sigmoid = 21'b111111111111100001010;
		14'b01001000011011:	sigmoid = 21'b111111111111100001010;
		14'b01001000011100:	sigmoid = 21'b111111111111100001010;
		14'b01001000011101:	sigmoid = 21'b111111111111100001011;
		14'b01001000011110:	sigmoid = 21'b111111111111100001011;
		14'b01001000011111:	sigmoid = 21'b111111111111100001100;
		14'b01001000100000:	sigmoid = 21'b111111111111100001100;
		14'b01001000100001:	sigmoid = 21'b111111111111100001101;
		14'b01001000100010:	sigmoid = 21'b111111111111100001101;
		14'b01001000100011:	sigmoid = 21'b111111111111100001110;
		14'b01001000100100:	sigmoid = 21'b111111111111100001110;
		14'b01001000100101:	sigmoid = 21'b111111111111100001111;
		14'b01001000100110:	sigmoid = 21'b111111111111100001111;
		14'b01001000100111:	sigmoid = 21'b111111111111100010000;
		14'b01001000101000:	sigmoid = 21'b111111111111100010000;
		14'b01001000101001:	sigmoid = 21'b111111111111100010001;
		14'b01001000101010:	sigmoid = 21'b111111111111100010001;
		14'b01001000101011:	sigmoid = 21'b111111111111100010010;
		14'b01001000101100:	sigmoid = 21'b111111111111100010010;
		14'b01001000101101:	sigmoid = 21'b111111111111100010010;
		14'b01001000101110:	sigmoid = 21'b111111111111100010011;
		14'b01001000101111:	sigmoid = 21'b111111111111100010011;
		14'b01001000110000:	sigmoid = 21'b111111111111100010100;
		14'b01001000110001:	sigmoid = 21'b111111111111100010100;
		14'b01001000110010:	sigmoid = 21'b111111111111100010101;
		14'b01001000110011:	sigmoid = 21'b111111111111100010101;
		14'b01001000110100:	sigmoid = 21'b111111111111100010110;
		14'b01001000110101:	sigmoid = 21'b111111111111100010110;
		14'b01001000110110:	sigmoid = 21'b111111111111100010111;
		14'b01001000110111:	sigmoid = 21'b111111111111100010111;
		14'b01001000111000:	sigmoid = 21'b111111111111100011000;
		14'b01001000111001:	sigmoid = 21'b111111111111100011000;
		14'b01001000111010:	sigmoid = 21'b111111111111100011000;
		14'b01001000111011:	sigmoid = 21'b111111111111100011001;
		14'b01001000111100:	sigmoid = 21'b111111111111100011001;
		14'b01001000111101:	sigmoid = 21'b111111111111100011010;
		14'b01001000111110:	sigmoid = 21'b111111111111100011010;
		14'b01001000111111:	sigmoid = 21'b111111111111100011011;
		14'b01001001000000:	sigmoid = 21'b111111111111100011011;
		14'b01001001000001:	sigmoid = 21'b111111111111100011100;
		14'b01001001000010:	sigmoid = 21'b111111111111100011100;
		14'b01001001000011:	sigmoid = 21'b111111111111100011100;
		14'b01001001000100:	sigmoid = 21'b111111111111100011101;
		14'b01001001000101:	sigmoid = 21'b111111111111100011101;
		14'b01001001000110:	sigmoid = 21'b111111111111100011110;
		14'b01001001000111:	sigmoid = 21'b111111111111100011110;
		14'b01001001001000:	sigmoid = 21'b111111111111100011111;
		14'b01001001001001:	sigmoid = 21'b111111111111100011111;
		14'b01001001001010:	sigmoid = 21'b111111111111100100000;
		14'b01001001001011:	sigmoid = 21'b111111111111100100000;
		14'b01001001001100:	sigmoid = 21'b111111111111100100000;
		14'b01001001001101:	sigmoid = 21'b111111111111100100001;
		14'b01001001001110:	sigmoid = 21'b111111111111100100001;
		14'b01001001001111:	sigmoid = 21'b111111111111100100010;
		14'b01001001010000:	sigmoid = 21'b111111111111100100010;
		14'b01001001010001:	sigmoid = 21'b111111111111100100011;
		14'b01001001010010:	sigmoid = 21'b111111111111100100011;
		14'b01001001010011:	sigmoid = 21'b111111111111100100011;
		14'b01001001010100:	sigmoid = 21'b111111111111100100100;
		14'b01001001010101:	sigmoid = 21'b111111111111100100100;
		14'b01001001010110:	sigmoid = 21'b111111111111100100101;
		14'b01001001010111:	sigmoid = 21'b111111111111100100101;
		14'b01001001011000:	sigmoid = 21'b111111111111100100110;
		14'b01001001011001:	sigmoid = 21'b111111111111100100110;
		14'b01001001011010:	sigmoid = 21'b111111111111100100110;
		14'b01001001011011:	sigmoid = 21'b111111111111100100111;
		14'b01001001011100:	sigmoid = 21'b111111111111100100111;
		14'b01001001011101:	sigmoid = 21'b111111111111100101000;
		14'b01001001011110:	sigmoid = 21'b111111111111100101000;
		14'b01001001011111:	sigmoid = 21'b111111111111100101001;
		14'b01001001100000:	sigmoid = 21'b111111111111100101001;
		14'b01001001100001:	sigmoid = 21'b111111111111100101001;
		14'b01001001100010:	sigmoid = 21'b111111111111100101010;
		14'b01001001100011:	sigmoid = 21'b111111111111100101010;
		14'b01001001100100:	sigmoid = 21'b111111111111100101011;
		14'b01001001100101:	sigmoid = 21'b111111111111100101011;
		14'b01001001100110:	sigmoid = 21'b111111111111100101011;
		14'b01001001100111:	sigmoid = 21'b111111111111100101100;
		14'b01001001101000:	sigmoid = 21'b111111111111100101100;
		14'b01001001101001:	sigmoid = 21'b111111111111100101101;
		14'b01001001101010:	sigmoid = 21'b111111111111100101101;
		14'b01001001101011:	sigmoid = 21'b111111111111100101110;
		14'b01001001101100:	sigmoid = 21'b111111111111100101110;
		14'b01001001101101:	sigmoid = 21'b111111111111100101110;
		14'b01001001101110:	sigmoid = 21'b111111111111100101111;
		14'b01001001101111:	sigmoid = 21'b111111111111100101111;
		14'b01001001110000:	sigmoid = 21'b111111111111100110000;
		14'b01001001110001:	sigmoid = 21'b111111111111100110000;
		14'b01001001110010:	sigmoid = 21'b111111111111100110000;
		14'b01001001110011:	sigmoid = 21'b111111111111100110001;
		14'b01001001110100:	sigmoid = 21'b111111111111100110001;
		14'b01001001110101:	sigmoid = 21'b111111111111100110010;
		14'b01001001110110:	sigmoid = 21'b111111111111100110010;
		14'b01001001110111:	sigmoid = 21'b111111111111100110010;
		14'b01001001111000:	sigmoid = 21'b111111111111100110011;
		14'b01001001111001:	sigmoid = 21'b111111111111100110011;
		14'b01001001111010:	sigmoid = 21'b111111111111100110100;
		14'b01001001111011:	sigmoid = 21'b111111111111100110100;
		14'b01001001111100:	sigmoid = 21'b111111111111100110100;
		14'b01001001111101:	sigmoid = 21'b111111111111100110101;
		14'b01001001111110:	sigmoid = 21'b111111111111100110101;
		14'b01001001111111:	sigmoid = 21'b111111111111100110110;
		14'b01001010000000:	sigmoid = 21'b111111111111100110110;
		14'b01001010000001:	sigmoid = 21'b111111111111100110110;
		14'b01001010000010:	sigmoid = 21'b111111111111100110111;
		14'b01001010000011:	sigmoid = 21'b111111111111100110111;
		14'b01001010000100:	sigmoid = 21'b111111111111100111000;
		14'b01001010000101:	sigmoid = 21'b111111111111100111000;
		14'b01001010000110:	sigmoid = 21'b111111111111100111000;
		14'b01001010000111:	sigmoid = 21'b111111111111100111001;
		14'b01001010001000:	sigmoid = 21'b111111111111100111001;
		14'b01001010001001:	sigmoid = 21'b111111111111100111001;
		14'b01001010001010:	sigmoid = 21'b111111111111100111010;
		14'b01001010001011:	sigmoid = 21'b111111111111100111010;
		14'b01001010001100:	sigmoid = 21'b111111111111100111011;
		14'b01001010001101:	sigmoid = 21'b111111111111100111011;
		14'b01001010001110:	sigmoid = 21'b111111111111100111011;
		14'b01001010001111:	sigmoid = 21'b111111111111100111100;
		14'b01001010010000:	sigmoid = 21'b111111111111100111100;
		14'b01001010010001:	sigmoid = 21'b111111111111100111101;
		14'b01001010010010:	sigmoid = 21'b111111111111100111101;
		14'b01001010010011:	sigmoid = 21'b111111111111100111101;
		14'b01001010010100:	sigmoid = 21'b111111111111100111110;
		14'b01001010010101:	sigmoid = 21'b111111111111100111110;
		14'b01001010010110:	sigmoid = 21'b111111111111100111110;
		14'b01001010010111:	sigmoid = 21'b111111111111100111111;
		14'b01001010011000:	sigmoid = 21'b111111111111100111111;
		14'b01001010011001:	sigmoid = 21'b111111111111101000000;
		14'b01001010011010:	sigmoid = 21'b111111111111101000000;
		14'b01001010011011:	sigmoid = 21'b111111111111101000000;
		14'b01001010011100:	sigmoid = 21'b111111111111101000001;
		14'b01001010011101:	sigmoid = 21'b111111111111101000001;
		14'b01001010011110:	sigmoid = 21'b111111111111101000001;
		14'b01001010011111:	sigmoid = 21'b111111111111101000010;
		14'b01001010100000:	sigmoid = 21'b111111111111101000010;
		14'b01001010100001:	sigmoid = 21'b111111111111101000011;
		14'b01001010100010:	sigmoid = 21'b111111111111101000011;
		14'b01001010100011:	sigmoid = 21'b111111111111101000011;
		14'b01001010100100:	sigmoid = 21'b111111111111101000100;
		14'b01001010100101:	sigmoid = 21'b111111111111101000100;
		14'b01001010100110:	sigmoid = 21'b111111111111101000100;
		14'b01001010100111:	sigmoid = 21'b111111111111101000101;
		14'b01001010101000:	sigmoid = 21'b111111111111101000101;
		14'b01001010101001:	sigmoid = 21'b111111111111101000101;
		14'b01001010101010:	sigmoid = 21'b111111111111101000110;
		14'b01001010101011:	sigmoid = 21'b111111111111101000110;
		14'b01001010101100:	sigmoid = 21'b111111111111101000111;
		14'b01001010101101:	sigmoid = 21'b111111111111101000111;
		14'b01001010101110:	sigmoid = 21'b111111111111101000111;
		14'b01001010101111:	sigmoid = 21'b111111111111101001000;
		14'b01001010110000:	sigmoid = 21'b111111111111101001000;
		14'b01001010110001:	sigmoid = 21'b111111111111101001000;
		14'b01001010110010:	sigmoid = 21'b111111111111101001001;
		14'b01001010110011:	sigmoid = 21'b111111111111101001001;
		14'b01001010110100:	sigmoid = 21'b111111111111101001001;
		14'b01001010110101:	sigmoid = 21'b111111111111101001010;
		14'b01001010110110:	sigmoid = 21'b111111111111101001010;
		14'b01001010110111:	sigmoid = 21'b111111111111101001010;
		14'b01001010111000:	sigmoid = 21'b111111111111101001011;
		14'b01001010111001:	sigmoid = 21'b111111111111101001011;
		14'b01001010111010:	sigmoid = 21'b111111111111101001100;
		14'b01001010111011:	sigmoid = 21'b111111111111101001100;
		14'b01001010111100:	sigmoid = 21'b111111111111101001100;
		14'b01001010111101:	sigmoid = 21'b111111111111101001101;
		14'b01001010111110:	sigmoid = 21'b111111111111101001101;
		14'b01001010111111:	sigmoid = 21'b111111111111101001101;
		14'b01001011000000:	sigmoid = 21'b111111111111101001110;
		14'b01001011000001:	sigmoid = 21'b111111111111101001110;
		14'b01001011000010:	sigmoid = 21'b111111111111101001110;
		14'b01001011000011:	sigmoid = 21'b111111111111101001111;
		14'b01001011000100:	sigmoid = 21'b111111111111101001111;
		14'b01001011000101:	sigmoid = 21'b111111111111101001111;
		14'b01001011000110:	sigmoid = 21'b111111111111101010000;
		14'b01001011000111:	sigmoid = 21'b111111111111101010000;
		14'b01001011001000:	sigmoid = 21'b111111111111101010000;
		14'b01001011001001:	sigmoid = 21'b111111111111101010001;
		14'b01001011001010:	sigmoid = 21'b111111111111101010001;
		14'b01001011001011:	sigmoid = 21'b111111111111101010001;
		14'b01001011001100:	sigmoid = 21'b111111111111101010010;
		14'b01001011001101:	sigmoid = 21'b111111111111101010010;
		14'b01001011001110:	sigmoid = 21'b111111111111101010010;
		14'b01001011001111:	sigmoid = 21'b111111111111101010011;
		14'b01001011010000:	sigmoid = 21'b111111111111101010011;
		14'b01001011010001:	sigmoid = 21'b111111111111101010011;
		14'b01001011010010:	sigmoid = 21'b111111111111101010100;
		14'b01001011010011:	sigmoid = 21'b111111111111101010100;
		14'b01001011010100:	sigmoid = 21'b111111111111101010100;
		14'b01001011010101:	sigmoid = 21'b111111111111101010101;
		14'b01001011010110:	sigmoid = 21'b111111111111101010101;
		14'b01001011010111:	sigmoid = 21'b111111111111101010101;
		14'b01001011011000:	sigmoid = 21'b111111111111101010110;
		14'b01001011011001:	sigmoid = 21'b111111111111101010110;
		14'b01001011011010:	sigmoid = 21'b111111111111101010110;
		14'b01001011011011:	sigmoid = 21'b111111111111101010111;
		14'b01001011011100:	sigmoid = 21'b111111111111101010111;
		14'b01001011011101:	sigmoid = 21'b111111111111101010111;
		14'b01001011011110:	sigmoid = 21'b111111111111101011000;
		14'b01001011011111:	sigmoid = 21'b111111111111101011000;
		14'b01001011100000:	sigmoid = 21'b111111111111101011000;
		14'b01001011100001:	sigmoid = 21'b111111111111101011001;
		14'b01001011100010:	sigmoid = 21'b111111111111101011001;
		14'b01001011100011:	sigmoid = 21'b111111111111101011001;
		14'b01001011100100:	sigmoid = 21'b111111111111101011010;
		14'b01001011100101:	sigmoid = 21'b111111111111101011010;
		14'b01001011100110:	sigmoid = 21'b111111111111101011010;
		14'b01001011100111:	sigmoid = 21'b111111111111101011011;
		14'b01001011101000:	sigmoid = 21'b111111111111101011011;
		14'b01001011101001:	sigmoid = 21'b111111111111101011011;
		14'b01001011101010:	sigmoid = 21'b111111111111101011100;
		14'b01001011101011:	sigmoid = 21'b111111111111101011100;
		14'b01001011101100:	sigmoid = 21'b111111111111101011100;
		14'b01001011101101:	sigmoid = 21'b111111111111101011101;
		14'b01001011101110:	sigmoid = 21'b111111111111101011101;
		14'b01001011101111:	sigmoid = 21'b111111111111101011101;
		14'b01001011110000:	sigmoid = 21'b111111111111101011110;
		14'b01001011110001:	sigmoid = 21'b111111111111101011110;
		14'b01001011110010:	sigmoid = 21'b111111111111101011110;
		14'b01001011110011:	sigmoid = 21'b111111111111101011110;
		14'b01001011110100:	sigmoid = 21'b111111111111101011111;
		14'b01001011110101:	sigmoid = 21'b111111111111101011111;
		14'b01001011110110:	sigmoid = 21'b111111111111101011111;
		14'b01001011110111:	sigmoid = 21'b111111111111101100000;
		14'b01001011111000:	sigmoid = 21'b111111111111101100000;
		14'b01001011111001:	sigmoid = 21'b111111111111101100000;
		14'b01001011111010:	sigmoid = 21'b111111111111101100001;
		14'b01001011111011:	sigmoid = 21'b111111111111101100001;
		14'b01001011111100:	sigmoid = 21'b111111111111101100001;
		14'b01001011111101:	sigmoid = 21'b111111111111101100010;
		14'b01001011111110:	sigmoid = 21'b111111111111101100010;
		14'b01001011111111:	sigmoid = 21'b111111111111101100010;
		14'b01001100000000:	sigmoid = 21'b111111111111101100011;
		14'b01001100000001:	sigmoid = 21'b111111111111101100011;
		14'b01001100000010:	sigmoid = 21'b111111111111101100011;
		14'b01001100000011:	sigmoid = 21'b111111111111101100011;
		14'b01001100000100:	sigmoid = 21'b111111111111101100100;
		14'b01001100000101:	sigmoid = 21'b111111111111101100100;
		14'b01001100000110:	sigmoid = 21'b111111111111101100100;
		14'b01001100000111:	sigmoid = 21'b111111111111101100101;
		14'b01001100001000:	sigmoid = 21'b111111111111101100101;
		14'b01001100001001:	sigmoid = 21'b111111111111101100101;
		14'b01001100001010:	sigmoid = 21'b111111111111101100110;
		14'b01001100001011:	sigmoid = 21'b111111111111101100110;
		14'b01001100001100:	sigmoid = 21'b111111111111101100110;
		14'b01001100001101:	sigmoid = 21'b111111111111101100110;
		14'b01001100001110:	sigmoid = 21'b111111111111101100111;
		14'b01001100001111:	sigmoid = 21'b111111111111101100111;
		14'b01001100010000:	sigmoid = 21'b111111111111101100111;
		14'b01001100010001:	sigmoid = 21'b111111111111101101000;
		14'b01001100010010:	sigmoid = 21'b111111111111101101000;
		14'b01001100010011:	sigmoid = 21'b111111111111101101000;
		14'b01001100010100:	sigmoid = 21'b111111111111101101001;
		14'b01001100010101:	sigmoid = 21'b111111111111101101001;
		14'b01001100010110:	sigmoid = 21'b111111111111101101001;
		14'b01001100010111:	sigmoid = 21'b111111111111101101001;
		14'b01001100011000:	sigmoid = 21'b111111111111101101010;
		14'b01001100011001:	sigmoid = 21'b111111111111101101010;
		14'b01001100011010:	sigmoid = 21'b111111111111101101010;
		14'b01001100011011:	sigmoid = 21'b111111111111101101011;
		14'b01001100011100:	sigmoid = 21'b111111111111101101011;
		14'b01001100011101:	sigmoid = 21'b111111111111101101011;
		14'b01001100011110:	sigmoid = 21'b111111111111101101011;
		14'b01001100011111:	sigmoid = 21'b111111111111101101100;
		14'b01001100100000:	sigmoid = 21'b111111111111101101100;
		14'b01001100100001:	sigmoid = 21'b111111111111101101100;
		14'b01001100100010:	sigmoid = 21'b111111111111101101101;
		14'b01001100100011:	sigmoid = 21'b111111111111101101101;
		14'b01001100100100:	sigmoid = 21'b111111111111101101101;
		14'b01001100100101:	sigmoid = 21'b111111111111101101101;
		14'b01001100100110:	sigmoid = 21'b111111111111101101110;
		14'b01001100100111:	sigmoid = 21'b111111111111101101110;
		14'b01001100101000:	sigmoid = 21'b111111111111101101110;
		14'b01001100101001:	sigmoid = 21'b111111111111101101111;
		14'b01001100101010:	sigmoid = 21'b111111111111101101111;
		14'b01001100101011:	sigmoid = 21'b111111111111101101111;
		14'b01001100101100:	sigmoid = 21'b111111111111101101111;
		14'b01001100101101:	sigmoid = 21'b111111111111101110000;
		14'b01001100101110:	sigmoid = 21'b111111111111101110000;
		14'b01001100101111:	sigmoid = 21'b111111111111101110000;
		14'b01001100110000:	sigmoid = 21'b111111111111101110001;
		14'b01001100110001:	sigmoid = 21'b111111111111101110001;
		14'b01001100110010:	sigmoid = 21'b111111111111101110001;
		14'b01001100110011:	sigmoid = 21'b111111111111101110001;
		14'b01001100110100:	sigmoid = 21'b111111111111101110010;
		14'b01001100110101:	sigmoid = 21'b111111111111101110010;
		14'b01001100110110:	sigmoid = 21'b111111111111101110010;
		14'b01001100110111:	sigmoid = 21'b111111111111101110011;
		14'b01001100111000:	sigmoid = 21'b111111111111101110011;
		14'b01001100111001:	sigmoid = 21'b111111111111101110011;
		14'b01001100111010:	sigmoid = 21'b111111111111101110011;
		14'b01001100111011:	sigmoid = 21'b111111111111101110100;
		14'b01001100111100:	sigmoid = 21'b111111111111101110100;
		14'b01001100111101:	sigmoid = 21'b111111111111101110100;
		14'b01001100111110:	sigmoid = 21'b111111111111101110100;
		14'b01001100111111:	sigmoid = 21'b111111111111101110101;
		14'b01001101000000:	sigmoid = 21'b111111111111101110101;
		14'b01001101000001:	sigmoid = 21'b111111111111101110101;
		14'b01001101000010:	sigmoid = 21'b111111111111101110110;
		14'b01001101000011:	sigmoid = 21'b111111111111101110110;
		14'b01001101000100:	sigmoid = 21'b111111111111101110110;
		14'b01001101000101:	sigmoid = 21'b111111111111101110110;
		14'b01001101000110:	sigmoid = 21'b111111111111101110111;
		14'b01001101000111:	sigmoid = 21'b111111111111101110111;
		14'b01001101001000:	sigmoid = 21'b111111111111101110111;
		14'b01001101001001:	sigmoid = 21'b111111111111101110111;
		14'b01001101001010:	sigmoid = 21'b111111111111101111000;
		14'b01001101001011:	sigmoid = 21'b111111111111101111000;
		14'b01001101001100:	sigmoid = 21'b111111111111101111000;
		14'b01001101001101:	sigmoid = 21'b111111111111101111000;
		14'b01001101001110:	sigmoid = 21'b111111111111101111001;
		14'b01001101001111:	sigmoid = 21'b111111111111101111001;
		14'b01001101010000:	sigmoid = 21'b111111111111101111001;
		14'b01001101010001:	sigmoid = 21'b111111111111101111010;
		14'b01001101010010:	sigmoid = 21'b111111111111101111010;
		14'b01001101010011:	sigmoid = 21'b111111111111101111010;
		14'b01001101010100:	sigmoid = 21'b111111111111101111010;
		14'b01001101010101:	sigmoid = 21'b111111111111101111011;
		14'b01001101010110:	sigmoid = 21'b111111111111101111011;
		14'b01001101010111:	sigmoid = 21'b111111111111101111011;
		14'b01001101011000:	sigmoid = 21'b111111111111101111011;
		14'b01001101011001:	sigmoid = 21'b111111111111101111100;
		14'b01001101011010:	sigmoid = 21'b111111111111101111100;
		14'b01001101011011:	sigmoid = 21'b111111111111101111100;
		14'b01001101011100:	sigmoid = 21'b111111111111101111100;
		14'b01001101011101:	sigmoid = 21'b111111111111101111101;
		14'b01001101011110:	sigmoid = 21'b111111111111101111101;
		14'b01001101011111:	sigmoid = 21'b111111111111101111101;
		14'b01001101100000:	sigmoid = 21'b111111111111101111101;
		14'b01001101100001:	sigmoid = 21'b111111111111101111110;
		14'b01001101100010:	sigmoid = 21'b111111111111101111110;
		14'b01001101100011:	sigmoid = 21'b111111111111101111110;
		14'b01001101100100:	sigmoid = 21'b111111111111101111110;
		14'b01001101100101:	sigmoid = 21'b111111111111101111111;
		14'b01001101100110:	sigmoid = 21'b111111111111101111111;
		14'b01001101100111:	sigmoid = 21'b111111111111101111111;
		14'b01001101101000:	sigmoid = 21'b111111111111101111111;
		14'b01001101101001:	sigmoid = 21'b111111111111110000000;
		14'b01001101101010:	sigmoid = 21'b111111111111110000000;
		14'b01001101101011:	sigmoid = 21'b111111111111110000000;
		14'b01001101101100:	sigmoid = 21'b111111111111110000000;
		14'b01001101101101:	sigmoid = 21'b111111111111110000001;
		14'b01001101101110:	sigmoid = 21'b111111111111110000001;
		14'b01001101101111:	sigmoid = 21'b111111111111110000001;
		14'b01001101110000:	sigmoid = 21'b111111111111110000001;
		14'b01001101110001:	sigmoid = 21'b111111111111110000010;
		14'b01001101110010:	sigmoid = 21'b111111111111110000010;
		14'b01001101110011:	sigmoid = 21'b111111111111110000010;
		14'b01001101110100:	sigmoid = 21'b111111111111110000010;
		14'b01001101110101:	sigmoid = 21'b111111111111110000011;
		14'b01001101110110:	sigmoid = 21'b111111111111110000011;
		14'b01001101110111:	sigmoid = 21'b111111111111110000011;
		14'b01001101111000:	sigmoid = 21'b111111111111110000011;
		14'b01001101111001:	sigmoid = 21'b111111111111110000100;
		14'b01001101111010:	sigmoid = 21'b111111111111110000100;
		14'b01001101111011:	sigmoid = 21'b111111111111110000100;
		14'b01001101111100:	sigmoid = 21'b111111111111110000100;
		14'b01001101111101:	sigmoid = 21'b111111111111110000101;
		14'b01001101111110:	sigmoid = 21'b111111111111110000101;
		14'b01001101111111:	sigmoid = 21'b111111111111110000101;
		14'b01001110000000:	sigmoid = 21'b111111111111110000101;
		14'b01001110000001:	sigmoid = 21'b111111111111110000101;
		14'b01001110000010:	sigmoid = 21'b111111111111110000110;
		14'b01001110000011:	sigmoid = 21'b111111111111110000110;
		14'b01001110000100:	sigmoid = 21'b111111111111110000110;
		14'b01001110000101:	sigmoid = 21'b111111111111110000110;
		14'b01001110000110:	sigmoid = 21'b111111111111110000111;
		14'b01001110000111:	sigmoid = 21'b111111111111110000111;
		14'b01001110001000:	sigmoid = 21'b111111111111110000111;
		14'b01001110001001:	sigmoid = 21'b111111111111110000111;
		14'b01001110001010:	sigmoid = 21'b111111111111110001000;
		14'b01001110001011:	sigmoid = 21'b111111111111110001000;
		14'b01001110001100:	sigmoid = 21'b111111111111110001000;
		14'b01001110001101:	sigmoid = 21'b111111111111110001000;
		14'b01001110001110:	sigmoid = 21'b111111111111110001001;
		14'b01001110001111:	sigmoid = 21'b111111111111110001001;
		14'b01001110010000:	sigmoid = 21'b111111111111110001001;
		14'b01001110010001:	sigmoid = 21'b111111111111110001001;
		14'b01001110010010:	sigmoid = 21'b111111111111110001001;
		14'b01001110010011:	sigmoid = 21'b111111111111110001010;
		14'b01001110010100:	sigmoid = 21'b111111111111110001010;
		14'b01001110010101:	sigmoid = 21'b111111111111110001010;
		14'b01001110010110:	sigmoid = 21'b111111111111110001010;
		14'b01001110010111:	sigmoid = 21'b111111111111110001011;
		14'b01001110011000:	sigmoid = 21'b111111111111110001011;
		14'b01001110011001:	sigmoid = 21'b111111111111110001011;
		14'b01001110011010:	sigmoid = 21'b111111111111110001011;
		14'b01001110011011:	sigmoid = 21'b111111111111110001100;
		14'b01001110011100:	sigmoid = 21'b111111111111110001100;
		14'b01001110011101:	sigmoid = 21'b111111111111110001100;
		14'b01001110011110:	sigmoid = 21'b111111111111110001100;
		14'b01001110011111:	sigmoid = 21'b111111111111110001100;
		14'b01001110100000:	sigmoid = 21'b111111111111110001101;
		14'b01001110100001:	sigmoid = 21'b111111111111110001101;
		14'b01001110100010:	sigmoid = 21'b111111111111110001101;
		14'b01001110100011:	sigmoid = 21'b111111111111110001101;
		14'b01001110100100:	sigmoid = 21'b111111111111110001110;
		14'b01001110100101:	sigmoid = 21'b111111111111110001110;
		14'b01001110100110:	sigmoid = 21'b111111111111110001110;
		14'b01001110100111:	sigmoid = 21'b111111111111110001110;
		14'b01001110101000:	sigmoid = 21'b111111111111110001110;
		14'b01001110101001:	sigmoid = 21'b111111111111110001111;
		14'b01001110101010:	sigmoid = 21'b111111111111110001111;
		14'b01001110101011:	sigmoid = 21'b111111111111110001111;
		14'b01001110101100:	sigmoid = 21'b111111111111110001111;
		14'b01001110101101:	sigmoid = 21'b111111111111110010000;
		14'b01001110101110:	sigmoid = 21'b111111111111110010000;
		14'b01001110101111:	sigmoid = 21'b111111111111110010000;
		14'b01001110110000:	sigmoid = 21'b111111111111110010000;
		14'b01001110110001:	sigmoid = 21'b111111111111110010000;
		14'b01001110110010:	sigmoid = 21'b111111111111110010001;
		14'b01001110110011:	sigmoid = 21'b111111111111110010001;
		14'b01001110110100:	sigmoid = 21'b111111111111110010001;
		14'b01001110110101:	sigmoid = 21'b111111111111110010001;
		14'b01001110110110:	sigmoid = 21'b111111111111110010001;
		14'b01001110110111:	sigmoid = 21'b111111111111110010010;
		14'b01001110111000:	sigmoid = 21'b111111111111110010010;
		14'b01001110111001:	sigmoid = 21'b111111111111110010010;
		14'b01001110111010:	sigmoid = 21'b111111111111110010010;
		14'b01001110111011:	sigmoid = 21'b111111111111110010011;
		14'b01001110111100:	sigmoid = 21'b111111111111110010011;
		14'b01001110111101:	sigmoid = 21'b111111111111110010011;
		14'b01001110111110:	sigmoid = 21'b111111111111110010011;
		14'b01001110111111:	sigmoid = 21'b111111111111110010011;
		14'b01001111000000:	sigmoid = 21'b111111111111110010100;
		14'b01001111000001:	sigmoid = 21'b111111111111110010100;
		14'b01001111000010:	sigmoid = 21'b111111111111110010100;
		14'b01001111000011:	sigmoid = 21'b111111111111110010100;
		14'b01001111000100:	sigmoid = 21'b111111111111110010100;
		14'b01001111000101:	sigmoid = 21'b111111111111110010101;
		14'b01001111000110:	sigmoid = 21'b111111111111110010101;
		14'b01001111000111:	sigmoid = 21'b111111111111110010101;
		14'b01001111001000:	sigmoid = 21'b111111111111110010101;
		14'b01001111001001:	sigmoid = 21'b111111111111110010101;
		14'b01001111001010:	sigmoid = 21'b111111111111110010110;
		14'b01001111001011:	sigmoid = 21'b111111111111110010110;
		14'b01001111001100:	sigmoid = 21'b111111111111110010110;
		14'b01001111001101:	sigmoid = 21'b111111111111110010110;
		14'b01001111001110:	sigmoid = 21'b111111111111110010111;
		14'b01001111001111:	sigmoid = 21'b111111111111110010111;
		14'b01001111010000:	sigmoid = 21'b111111111111110010111;
		14'b01001111010001:	sigmoid = 21'b111111111111110010111;
		14'b01001111010010:	sigmoid = 21'b111111111111110010111;
		14'b01001111010011:	sigmoid = 21'b111111111111110011000;
		14'b01001111010100:	sigmoid = 21'b111111111111110011000;
		14'b01001111010101:	sigmoid = 21'b111111111111110011000;
		14'b01001111010110:	sigmoid = 21'b111111111111110011000;
		14'b01001111010111:	sigmoid = 21'b111111111111110011000;
		14'b01001111011000:	sigmoid = 21'b111111111111110011001;
		14'b01001111011001:	sigmoid = 21'b111111111111110011001;
		14'b01001111011010:	sigmoid = 21'b111111111111110011001;
		14'b01001111011011:	sigmoid = 21'b111111111111110011001;
		14'b01001111011100:	sigmoid = 21'b111111111111110011001;
		14'b01001111011101:	sigmoid = 21'b111111111111110011010;
		14'b01001111011110:	sigmoid = 21'b111111111111110011010;
		14'b01001111011111:	sigmoid = 21'b111111111111110011010;
		14'b01001111100000:	sigmoid = 21'b111111111111110011010;
		14'b01001111100001:	sigmoid = 21'b111111111111110011010;
		14'b01001111100010:	sigmoid = 21'b111111111111110011011;
		14'b01001111100011:	sigmoid = 21'b111111111111110011011;
		14'b01001111100100:	sigmoid = 21'b111111111111110011011;
		14'b01001111100101:	sigmoid = 21'b111111111111110011011;
		14'b01001111100110:	sigmoid = 21'b111111111111110011011;
		14'b01001111100111:	sigmoid = 21'b111111111111110011100;
		14'b01001111101000:	sigmoid = 21'b111111111111110011100;
		14'b01001111101001:	sigmoid = 21'b111111111111110011100;
		14'b01001111101010:	sigmoid = 21'b111111111111110011100;
		14'b01001111101011:	sigmoid = 21'b111111111111110011100;
		14'b01001111101100:	sigmoid = 21'b111111111111110011101;
		14'b01001111101101:	sigmoid = 21'b111111111111110011101;
		14'b01001111101110:	sigmoid = 21'b111111111111110011101;
		14'b01001111101111:	sigmoid = 21'b111111111111110011101;
		14'b01001111110000:	sigmoid = 21'b111111111111110011101;
		14'b01001111110001:	sigmoid = 21'b111111111111110011101;
		14'b01001111110010:	sigmoid = 21'b111111111111110011110;
		14'b01001111110011:	sigmoid = 21'b111111111111110011110;
		14'b01001111110100:	sigmoid = 21'b111111111111110011110;
		14'b01001111110101:	sigmoid = 21'b111111111111110011110;
		14'b01001111110110:	sigmoid = 21'b111111111111110011110;
		14'b01001111110111:	sigmoid = 21'b111111111111110011111;
		14'b01001111111000:	sigmoid = 21'b111111111111110011111;
		14'b01001111111001:	sigmoid = 21'b111111111111110011111;
		14'b01001111111010:	sigmoid = 21'b111111111111110011111;
		14'b01001111111011:	sigmoid = 21'b111111111111110011111;
		14'b01001111111100:	sigmoid = 21'b111111111111110100000;
		14'b01001111111101:	sigmoid = 21'b111111111111110100000;
		14'b01001111111110:	sigmoid = 21'b111111111111110100000;
		14'b01001111111111:	sigmoid = 21'b111111111111110100000;
		14'b01010000000000:	sigmoid = 21'b111111111111110100000;
		14'b01010000000001:	sigmoid = 21'b111111111111110100000;
		14'b01010000000010:	sigmoid = 21'b111111111111110100001;
		14'b01010000000011:	sigmoid = 21'b111111111111110100001;
		14'b01010000000100:	sigmoid = 21'b111111111111110100001;
		14'b01010000000101:	sigmoid = 21'b111111111111110100001;
		14'b01010000000110:	sigmoid = 21'b111111111111110100001;
		14'b01010000000111:	sigmoid = 21'b111111111111110100010;
		14'b01010000001000:	sigmoid = 21'b111111111111110100010;
		14'b01010000001001:	sigmoid = 21'b111111111111110100010;
		14'b01010000001010:	sigmoid = 21'b111111111111110100010;
		14'b01010000001011:	sigmoid = 21'b111111111111110100010;
		14'b01010000001100:	sigmoid = 21'b111111111111110100010;
		14'b01010000001101:	sigmoid = 21'b111111111111110100011;
		14'b01010000001110:	sigmoid = 21'b111111111111110100011;
		14'b01010000001111:	sigmoid = 21'b111111111111110100011;
		14'b01010000010000:	sigmoid = 21'b111111111111110100011;
		14'b01010000010001:	sigmoid = 21'b111111111111110100011;
		14'b01010000010010:	sigmoid = 21'b111111111111110100100;
		14'b01010000010011:	sigmoid = 21'b111111111111110100100;
		14'b01010000010100:	sigmoid = 21'b111111111111110100100;
		14'b01010000010101:	sigmoid = 21'b111111111111110100100;
		14'b01010000010110:	sigmoid = 21'b111111111111110100100;
		14'b01010000010111:	sigmoid = 21'b111111111111110100100;
		14'b01010000011000:	sigmoid = 21'b111111111111110100101;
		14'b01010000011001:	sigmoid = 21'b111111111111110100101;
		14'b01010000011010:	sigmoid = 21'b111111111111110100101;
		14'b01010000011011:	sigmoid = 21'b111111111111110100101;
		14'b01010000011100:	sigmoid = 21'b111111111111110100101;
		14'b01010000011101:	sigmoid = 21'b111111111111110100110;
		14'b01010000011110:	sigmoid = 21'b111111111111110100110;
		14'b01010000011111:	sigmoid = 21'b111111111111110100110;
		14'b01010000100000:	sigmoid = 21'b111111111111110100110;
		14'b01010000100001:	sigmoid = 21'b111111111111110100110;
		14'b01010000100010:	sigmoid = 21'b111111111111110100110;
		14'b01010000100011:	sigmoid = 21'b111111111111110100111;
		14'b01010000100100:	sigmoid = 21'b111111111111110100111;
		14'b01010000100101:	sigmoid = 21'b111111111111110100111;
		14'b01010000100110:	sigmoid = 21'b111111111111110100111;
		14'b01010000100111:	sigmoid = 21'b111111111111110100111;
		14'b01010000101000:	sigmoid = 21'b111111111111110100111;
		14'b01010000101001:	sigmoid = 21'b111111111111110101000;
		14'b01010000101010:	sigmoid = 21'b111111111111110101000;
		14'b01010000101011:	sigmoid = 21'b111111111111110101000;
		14'b01010000101100:	sigmoid = 21'b111111111111110101000;
		14'b01010000101101:	sigmoid = 21'b111111111111110101000;
		14'b01010000101110:	sigmoid = 21'b111111111111110101000;
		14'b01010000101111:	sigmoid = 21'b111111111111110101001;
		14'b01010000110000:	sigmoid = 21'b111111111111110101001;
		14'b01010000110001:	sigmoid = 21'b111111111111110101001;
		14'b01010000110010:	sigmoid = 21'b111111111111110101001;
		14'b01010000110011:	sigmoid = 21'b111111111111110101001;
		14'b01010000110100:	sigmoid = 21'b111111111111110101001;
		14'b01010000110101:	sigmoid = 21'b111111111111110101010;
		14'b01010000110110:	sigmoid = 21'b111111111111110101010;
		14'b01010000110111:	sigmoid = 21'b111111111111110101010;
		14'b01010000111000:	sigmoid = 21'b111111111111110101010;
		14'b01010000111001:	sigmoid = 21'b111111111111110101010;
		14'b01010000111010:	sigmoid = 21'b111111111111110101010;
		14'b01010000111011:	sigmoid = 21'b111111111111110101011;
		14'b01010000111100:	sigmoid = 21'b111111111111110101011;
		14'b01010000111101:	sigmoid = 21'b111111111111110101011;
		14'b01010000111110:	sigmoid = 21'b111111111111110101011;
		14'b01010000111111:	sigmoid = 21'b111111111111110101011;
		14'b01010001000000:	sigmoid = 21'b111111111111110101011;
		14'b01010001000001:	sigmoid = 21'b111111111111110101100;
		14'b01010001000010:	sigmoid = 21'b111111111111110101100;
		14'b01010001000011:	sigmoid = 21'b111111111111110101100;
		14'b01010001000100:	sigmoid = 21'b111111111111110101100;
		14'b01010001000101:	sigmoid = 21'b111111111111110101100;
		14'b01010001000110:	sigmoid = 21'b111111111111110101100;
		14'b01010001000111:	sigmoid = 21'b111111111111110101101;
		14'b01010001001000:	sigmoid = 21'b111111111111110101101;
		14'b01010001001001:	sigmoid = 21'b111111111111110101101;
		14'b01010001001010:	sigmoid = 21'b111111111111110101101;
		14'b01010001001011:	sigmoid = 21'b111111111111110101101;
		14'b01010001001100:	sigmoid = 21'b111111111111110101101;
		14'b01010001001101:	sigmoid = 21'b111111111111110101110;
		14'b01010001001110:	sigmoid = 21'b111111111111110101110;
		14'b01010001001111:	sigmoid = 21'b111111111111110101110;
		14'b01010001010000:	sigmoid = 21'b111111111111110101110;
		14'b01010001010001:	sigmoid = 21'b111111111111110101110;
		14'b01010001010010:	sigmoid = 21'b111111111111110101110;
		14'b01010001010011:	sigmoid = 21'b111111111111110101111;
		14'b01010001010100:	sigmoid = 21'b111111111111110101111;
		14'b01010001010101:	sigmoid = 21'b111111111111110101111;
		14'b01010001010110:	sigmoid = 21'b111111111111110101111;
		14'b01010001010111:	sigmoid = 21'b111111111111110101111;
		14'b01010001011000:	sigmoid = 21'b111111111111110101111;
		14'b01010001011001:	sigmoid = 21'b111111111111110101111;
		14'b01010001011010:	sigmoid = 21'b111111111111110110000;
		14'b01010001011011:	sigmoid = 21'b111111111111110110000;
		14'b01010001011100:	sigmoid = 21'b111111111111110110000;
		14'b01010001011101:	sigmoid = 21'b111111111111110110000;
		14'b01010001011110:	sigmoid = 21'b111111111111110110000;
		14'b01010001011111:	sigmoid = 21'b111111111111110110000;
		14'b01010001100000:	sigmoid = 21'b111111111111110110001;
		14'b01010001100001:	sigmoid = 21'b111111111111110110001;
		14'b01010001100010:	sigmoid = 21'b111111111111110110001;
		14'b01010001100011:	sigmoid = 21'b111111111111110110001;
		14'b01010001100100:	sigmoid = 21'b111111111111110110001;
		14'b01010001100101:	sigmoid = 21'b111111111111110110001;
		14'b01010001100110:	sigmoid = 21'b111111111111110110001;
		14'b01010001100111:	sigmoid = 21'b111111111111110110010;
		14'b01010001101000:	sigmoid = 21'b111111111111110110010;
		14'b01010001101001:	sigmoid = 21'b111111111111110110010;
		14'b01010001101010:	sigmoid = 21'b111111111111110110010;
		14'b01010001101011:	sigmoid = 21'b111111111111110110010;
		14'b01010001101100:	sigmoid = 21'b111111111111110110010;
		14'b01010001101101:	sigmoid = 21'b111111111111110110011;
		14'b01010001101110:	sigmoid = 21'b111111111111110110011;
		14'b01010001101111:	sigmoid = 21'b111111111111110110011;
		14'b01010001110000:	sigmoid = 21'b111111111111110110011;
		14'b01010001110001:	sigmoid = 21'b111111111111110110011;
		14'b01010001110010:	sigmoid = 21'b111111111111110110011;
		14'b01010001110011:	sigmoid = 21'b111111111111110110011;
		14'b01010001110100:	sigmoid = 21'b111111111111110110100;
		14'b01010001110101:	sigmoid = 21'b111111111111110110100;
		14'b01010001110110:	sigmoid = 21'b111111111111110110100;
		14'b01010001110111:	sigmoid = 21'b111111111111110110100;
		14'b01010001111000:	sigmoid = 21'b111111111111110110100;
		14'b01010001111001:	sigmoid = 21'b111111111111110110100;
		14'b01010001111010:	sigmoid = 21'b111111111111110110100;
		14'b01010001111011:	sigmoid = 21'b111111111111110110101;
		14'b01010001111100:	sigmoid = 21'b111111111111110110101;
		14'b01010001111101:	sigmoid = 21'b111111111111110110101;
		14'b01010001111110:	sigmoid = 21'b111111111111110110101;
		14'b01010001111111:	sigmoid = 21'b111111111111110110101;
		14'b01010010000000:	sigmoid = 21'b111111111111110110101;
		14'b01010010000001:	sigmoid = 21'b111111111111110110101;
		14'b01010010000010:	sigmoid = 21'b111111111111110110110;
		14'b01010010000011:	sigmoid = 21'b111111111111110110110;
		14'b01010010000100:	sigmoid = 21'b111111111111110110110;
		14'b01010010000101:	sigmoid = 21'b111111111111110110110;
		14'b01010010000110:	sigmoid = 21'b111111111111110110110;
		14'b01010010000111:	sigmoid = 21'b111111111111110110110;
		14'b01010010001000:	sigmoid = 21'b111111111111110110111;
		14'b01010010001001:	sigmoid = 21'b111111111111110110111;
		14'b01010010001010:	sigmoid = 21'b111111111111110110111;
		14'b01010010001011:	sigmoid = 21'b111111111111110110111;
		14'b01010010001100:	sigmoid = 21'b111111111111110110111;
		14'b01010010001101:	sigmoid = 21'b111111111111110110111;
		14'b01010010001110:	sigmoid = 21'b111111111111110110111;
		14'b01010010001111:	sigmoid = 21'b111111111111110110111;
		14'b01010010010000:	sigmoid = 21'b111111111111110111000;
		14'b01010010010001:	sigmoid = 21'b111111111111110111000;
		14'b01010010010010:	sigmoid = 21'b111111111111110111000;
		14'b01010010010011:	sigmoid = 21'b111111111111110111000;
		14'b01010010010100:	sigmoid = 21'b111111111111110111000;
		14'b01010010010101:	sigmoid = 21'b111111111111110111000;
		14'b01010010010110:	sigmoid = 21'b111111111111110111000;
		14'b01010010010111:	sigmoid = 21'b111111111111110111001;
		14'b01010010011000:	sigmoid = 21'b111111111111110111001;
		14'b01010010011001:	sigmoid = 21'b111111111111110111001;
		14'b01010010011010:	sigmoid = 21'b111111111111110111001;
		14'b01010010011011:	sigmoid = 21'b111111111111110111001;
		14'b01010010011100:	sigmoid = 21'b111111111111110111001;
		14'b01010010011101:	sigmoid = 21'b111111111111110111001;
		14'b01010010011110:	sigmoid = 21'b111111111111110111010;
		14'b01010010011111:	sigmoid = 21'b111111111111110111010;
		14'b01010010100000:	sigmoid = 21'b111111111111110111010;
		14'b01010010100001:	sigmoid = 21'b111111111111110111010;
		14'b01010010100010:	sigmoid = 21'b111111111111110111010;
		14'b01010010100011:	sigmoid = 21'b111111111111110111010;
		14'b01010010100100:	sigmoid = 21'b111111111111110111010;
		14'b01010010100101:	sigmoid = 21'b111111111111110111011;
		14'b01010010100110:	sigmoid = 21'b111111111111110111011;
		14'b01010010100111:	sigmoid = 21'b111111111111110111011;
		14'b01010010101000:	sigmoid = 21'b111111111111110111011;
		14'b01010010101001:	sigmoid = 21'b111111111111110111011;
		14'b01010010101010:	sigmoid = 21'b111111111111110111011;
		14'b01010010101011:	sigmoid = 21'b111111111111110111011;
		14'b01010010101100:	sigmoid = 21'b111111111111110111011;
		14'b01010010101101:	sigmoid = 21'b111111111111110111100;
		14'b01010010101110:	sigmoid = 21'b111111111111110111100;
		14'b01010010101111:	sigmoid = 21'b111111111111110111100;
		14'b01010010110000:	sigmoid = 21'b111111111111110111100;
		14'b01010010110001:	sigmoid = 21'b111111111111110111100;
		14'b01010010110010:	sigmoid = 21'b111111111111110111100;
		14'b01010010110011:	sigmoid = 21'b111111111111110111100;
		14'b01010010110100:	sigmoid = 21'b111111111111110111101;
		14'b01010010110101:	sigmoid = 21'b111111111111110111101;
		14'b01010010110110:	sigmoid = 21'b111111111111110111101;
		14'b01010010110111:	sigmoid = 21'b111111111111110111101;
		14'b01010010111000:	sigmoid = 21'b111111111111110111101;
		14'b01010010111001:	sigmoid = 21'b111111111111110111101;
		14'b01010010111010:	sigmoid = 21'b111111111111110111101;
		14'b01010010111011:	sigmoid = 21'b111111111111110111101;
		14'b01010010111100:	sigmoid = 21'b111111111111110111110;
		14'b01010010111101:	sigmoid = 21'b111111111111110111110;
		14'b01010010111110:	sigmoid = 21'b111111111111110111110;
		14'b01010010111111:	sigmoid = 21'b111111111111110111110;
		14'b01010011000000:	sigmoid = 21'b111111111111110111110;
		14'b01010011000001:	sigmoid = 21'b111111111111110111110;
		14'b01010011000010:	sigmoid = 21'b111111111111110111110;
		14'b01010011000011:	sigmoid = 21'b111111111111110111110;
		14'b01010011000100:	sigmoid = 21'b111111111111110111111;
		14'b01010011000101:	sigmoid = 21'b111111111111110111111;
		14'b01010011000110:	sigmoid = 21'b111111111111110111111;
		14'b01010011000111:	sigmoid = 21'b111111111111110111111;
		14'b01010011001000:	sigmoid = 21'b111111111111110111111;
		14'b01010011001001:	sigmoid = 21'b111111111111110111111;
		14'b01010011001010:	sigmoid = 21'b111111111111110111111;
		14'b01010011001011:	sigmoid = 21'b111111111111110111111;
		14'b01010011001100:	sigmoid = 21'b111111111111111000000;
		14'b01010011001101:	sigmoid = 21'b111111111111111000000;
		14'b01010011001110:	sigmoid = 21'b111111111111111000000;
		14'b01010011001111:	sigmoid = 21'b111111111111111000000;
		14'b01010011010000:	sigmoid = 21'b111111111111111000000;
		14'b01010011010001:	sigmoid = 21'b111111111111111000000;
		14'b01010011010010:	sigmoid = 21'b111111111111111000000;
		14'b01010011010011:	sigmoid = 21'b111111111111111000000;
		14'b01010011010100:	sigmoid = 21'b111111111111111000001;
		14'b01010011010101:	sigmoid = 21'b111111111111111000001;
		14'b01010011010110:	sigmoid = 21'b111111111111111000001;
		14'b01010011010111:	sigmoid = 21'b111111111111111000001;
		14'b01010011011000:	sigmoid = 21'b111111111111111000001;
		14'b01010011011001:	sigmoid = 21'b111111111111111000001;
		14'b01010011011010:	sigmoid = 21'b111111111111111000001;
		14'b01010011011011:	sigmoid = 21'b111111111111111000001;
		14'b01010011011100:	sigmoid = 21'b111111111111111000010;
		14'b01010011011101:	sigmoid = 21'b111111111111111000010;
		14'b01010011011110:	sigmoid = 21'b111111111111111000010;
		14'b01010011011111:	sigmoid = 21'b111111111111111000010;
		14'b01010011100000:	sigmoid = 21'b111111111111111000010;
		14'b01010011100001:	sigmoid = 21'b111111111111111000010;
		14'b01010011100010:	sigmoid = 21'b111111111111111000010;
		14'b01010011100011:	sigmoid = 21'b111111111111111000010;
		14'b01010011100100:	sigmoid = 21'b111111111111111000011;
		14'b01010011100101:	sigmoid = 21'b111111111111111000011;
		14'b01010011100110:	sigmoid = 21'b111111111111111000011;
		14'b01010011100111:	sigmoid = 21'b111111111111111000011;
		14'b01010011101000:	sigmoid = 21'b111111111111111000011;
		14'b01010011101001:	sigmoid = 21'b111111111111111000011;
		14'b01010011101010:	sigmoid = 21'b111111111111111000011;
		14'b01010011101011:	sigmoid = 21'b111111111111111000011;
		14'b01010011101100:	sigmoid = 21'b111111111111111000011;
		14'b01010011101101:	sigmoid = 21'b111111111111111000100;
		14'b01010011101110:	sigmoid = 21'b111111111111111000100;
		14'b01010011101111:	sigmoid = 21'b111111111111111000100;
		14'b01010011110000:	sigmoid = 21'b111111111111111000100;
		14'b01010011110001:	sigmoid = 21'b111111111111111000100;
		14'b01010011110010:	sigmoid = 21'b111111111111111000100;
		14'b01010011110011:	sigmoid = 21'b111111111111111000100;
		14'b01010011110100:	sigmoid = 21'b111111111111111000100;
		14'b01010011110101:	sigmoid = 21'b111111111111111000100;
		14'b01010011110110:	sigmoid = 21'b111111111111111000101;
		14'b01010011110111:	sigmoid = 21'b111111111111111000101;
		14'b01010011111000:	sigmoid = 21'b111111111111111000101;
		14'b01010011111001:	sigmoid = 21'b111111111111111000101;
		14'b01010011111010:	sigmoid = 21'b111111111111111000101;
		14'b01010011111011:	sigmoid = 21'b111111111111111000101;
		14'b01010011111100:	sigmoid = 21'b111111111111111000101;
		14'b01010011111101:	sigmoid = 21'b111111111111111000101;
		14'b01010011111110:	sigmoid = 21'b111111111111111000110;
		14'b01010011111111:	sigmoid = 21'b111111111111111000110;
		14'b01010100000000:	sigmoid = 21'b111111111111111000110;
		14'b01010100000001:	sigmoid = 21'b111111111111111000110;
		14'b01010100000010:	sigmoid = 21'b111111111111111000110;
		14'b01010100000011:	sigmoid = 21'b111111111111111000110;
		14'b01010100000100:	sigmoid = 21'b111111111111111000110;
		14'b01010100000101:	sigmoid = 21'b111111111111111000110;
		14'b01010100000110:	sigmoid = 21'b111111111111111000110;
		14'b01010100000111:	sigmoid = 21'b111111111111111000111;
		14'b01010100001000:	sigmoid = 21'b111111111111111000111;
		14'b01010100001001:	sigmoid = 21'b111111111111111000111;
		14'b01010100001010:	sigmoid = 21'b111111111111111000111;
		14'b01010100001011:	sigmoid = 21'b111111111111111000111;
		14'b01010100001100:	sigmoid = 21'b111111111111111000111;
		14'b01010100001101:	sigmoid = 21'b111111111111111000111;
		14'b01010100001110:	sigmoid = 21'b111111111111111000111;
		14'b01010100001111:	sigmoid = 21'b111111111111111000111;
		14'b01010100010000:	sigmoid = 21'b111111111111111001000;
		14'b01010100010001:	sigmoid = 21'b111111111111111001000;
		14'b01010100010010:	sigmoid = 21'b111111111111111001000;
		14'b01010100010011:	sigmoid = 21'b111111111111111001000;
		14'b01010100010100:	sigmoid = 21'b111111111111111001000;
		14'b01010100010101:	sigmoid = 21'b111111111111111001000;
		14'b01010100010110:	sigmoid = 21'b111111111111111001000;
		14'b01010100010111:	sigmoid = 21'b111111111111111001000;
		14'b01010100011000:	sigmoid = 21'b111111111111111001000;
		14'b01010100011001:	sigmoid = 21'b111111111111111001001;
		14'b01010100011010:	sigmoid = 21'b111111111111111001001;
		14'b01010100011011:	sigmoid = 21'b111111111111111001001;
		14'b01010100011100:	sigmoid = 21'b111111111111111001001;
		14'b01010100011101:	sigmoid = 21'b111111111111111001001;
		14'b01010100011110:	sigmoid = 21'b111111111111111001001;
		14'b01010100011111:	sigmoid = 21'b111111111111111001001;
		14'b01010100100000:	sigmoid = 21'b111111111111111001001;
		14'b01010100100001:	sigmoid = 21'b111111111111111001001;
		14'b01010100100010:	sigmoid = 21'b111111111111111001001;
		14'b01010100100011:	sigmoid = 21'b111111111111111001010;
		14'b01010100100100:	sigmoid = 21'b111111111111111001010;
		14'b01010100100101:	sigmoid = 21'b111111111111111001010;
		14'b01010100100110:	sigmoid = 21'b111111111111111001010;
		14'b01010100100111:	sigmoid = 21'b111111111111111001010;
		14'b01010100101000:	sigmoid = 21'b111111111111111001010;
		14'b01010100101001:	sigmoid = 21'b111111111111111001010;
		14'b01010100101010:	sigmoid = 21'b111111111111111001010;
		14'b01010100101011:	sigmoid = 21'b111111111111111001010;
		14'b01010100101100:	sigmoid = 21'b111111111111111001011;
		14'b01010100101101:	sigmoid = 21'b111111111111111001011;
		14'b01010100101110:	sigmoid = 21'b111111111111111001011;
		14'b01010100101111:	sigmoid = 21'b111111111111111001011;
		14'b01010100110000:	sigmoid = 21'b111111111111111001011;
		14'b01010100110001:	sigmoid = 21'b111111111111111001011;
		14'b01010100110010:	sigmoid = 21'b111111111111111001011;
		14'b01010100110011:	sigmoid = 21'b111111111111111001011;
		14'b01010100110100:	sigmoid = 21'b111111111111111001011;
		14'b01010100110101:	sigmoid = 21'b111111111111111001011;
		14'b01010100110110:	sigmoid = 21'b111111111111111001100;
		14'b01010100110111:	sigmoid = 21'b111111111111111001100;
		14'b01010100111000:	sigmoid = 21'b111111111111111001100;
		14'b01010100111001:	sigmoid = 21'b111111111111111001100;
		14'b01010100111010:	sigmoid = 21'b111111111111111001100;
		14'b01010100111011:	sigmoid = 21'b111111111111111001100;
		14'b01010100111100:	sigmoid = 21'b111111111111111001100;
		14'b01010100111101:	sigmoid = 21'b111111111111111001100;
		14'b01010100111110:	sigmoid = 21'b111111111111111001100;
		14'b01010100111111:	sigmoid = 21'b111111111111111001100;
		14'b01010101000000:	sigmoid = 21'b111111111111111001101;
		14'b01010101000001:	sigmoid = 21'b111111111111111001101;
		14'b01010101000010:	sigmoid = 21'b111111111111111001101;
		14'b01010101000011:	sigmoid = 21'b111111111111111001101;
		14'b01010101000100:	sigmoid = 21'b111111111111111001101;
		14'b01010101000101:	sigmoid = 21'b111111111111111001101;
		14'b01010101000110:	sigmoid = 21'b111111111111111001101;
		14'b01010101000111:	sigmoid = 21'b111111111111111001101;
		14'b01010101001000:	sigmoid = 21'b111111111111111001101;
		14'b01010101001001:	sigmoid = 21'b111111111111111001101;
		14'b01010101001010:	sigmoid = 21'b111111111111111001110;
		14'b01010101001011:	sigmoid = 21'b111111111111111001110;
		14'b01010101001100:	sigmoid = 21'b111111111111111001110;
		14'b01010101001101:	sigmoid = 21'b111111111111111001110;
		14'b01010101001110:	sigmoid = 21'b111111111111111001110;
		14'b01010101001111:	sigmoid = 21'b111111111111111001110;
		14'b01010101010000:	sigmoid = 21'b111111111111111001110;
		14'b01010101010001:	sigmoid = 21'b111111111111111001110;
		14'b01010101010010:	sigmoid = 21'b111111111111111001110;
		14'b01010101010011:	sigmoid = 21'b111111111111111001110;
		14'b01010101010100:	sigmoid = 21'b111111111111111001110;
		14'b01010101010101:	sigmoid = 21'b111111111111111001111;
		14'b01010101010110:	sigmoid = 21'b111111111111111001111;
		14'b01010101010111:	sigmoid = 21'b111111111111111001111;
		14'b01010101011000:	sigmoid = 21'b111111111111111001111;
		14'b01010101011001:	sigmoid = 21'b111111111111111001111;
		14'b01010101011010:	sigmoid = 21'b111111111111111001111;
		14'b01010101011011:	sigmoid = 21'b111111111111111001111;
		14'b01010101011100:	sigmoid = 21'b111111111111111001111;
		14'b01010101011101:	sigmoid = 21'b111111111111111001111;
		14'b01010101011110:	sigmoid = 21'b111111111111111001111;
		14'b01010101011111:	sigmoid = 21'b111111111111111010000;
		14'b01010101100000:	sigmoid = 21'b111111111111111010000;
		14'b01010101100001:	sigmoid = 21'b111111111111111010000;
		14'b01010101100010:	sigmoid = 21'b111111111111111010000;
		14'b01010101100011:	sigmoid = 21'b111111111111111010000;
		14'b01010101100100:	sigmoid = 21'b111111111111111010000;
		14'b01010101100101:	sigmoid = 21'b111111111111111010000;
		14'b01010101100110:	sigmoid = 21'b111111111111111010000;
		14'b01010101100111:	sigmoid = 21'b111111111111111010000;
		14'b01010101101000:	sigmoid = 21'b111111111111111010000;
		14'b01010101101001:	sigmoid = 21'b111111111111111010000;
		14'b01010101101010:	sigmoid = 21'b111111111111111010001;
		14'b01010101101011:	sigmoid = 21'b111111111111111010001;
		14'b01010101101100:	sigmoid = 21'b111111111111111010001;
		14'b01010101101101:	sigmoid = 21'b111111111111111010001;
		14'b01010101101110:	sigmoid = 21'b111111111111111010001;
		14'b01010101101111:	sigmoid = 21'b111111111111111010001;
		14'b01010101110000:	sigmoid = 21'b111111111111111010001;
		14'b01010101110001:	sigmoid = 21'b111111111111111010001;
		14'b01010101110010:	sigmoid = 21'b111111111111111010001;
		14'b01010101110011:	sigmoid = 21'b111111111111111010001;
		14'b01010101110100:	sigmoid = 21'b111111111111111010001;
		14'b01010101110101:	sigmoid = 21'b111111111111111010010;
		14'b01010101110110:	sigmoid = 21'b111111111111111010010;
		14'b01010101110111:	sigmoid = 21'b111111111111111010010;
		14'b01010101111000:	sigmoid = 21'b111111111111111010010;
		14'b01010101111001:	sigmoid = 21'b111111111111111010010;
		14'b01010101111010:	sigmoid = 21'b111111111111111010010;
		14'b01010101111011:	sigmoid = 21'b111111111111111010010;
		14'b01010101111100:	sigmoid = 21'b111111111111111010010;
		14'b01010101111101:	sigmoid = 21'b111111111111111010010;
		14'b01010101111110:	sigmoid = 21'b111111111111111010010;
		14'b01010101111111:	sigmoid = 21'b111111111111111010010;
		14'b01010110000000:	sigmoid = 21'b111111111111111010011;
		14'b01010110000001:	sigmoid = 21'b111111111111111010011;
		14'b01010110000010:	sigmoid = 21'b111111111111111010011;
		14'b01010110000011:	sigmoid = 21'b111111111111111010011;
		14'b01010110000100:	sigmoid = 21'b111111111111111010011;
		14'b01010110000101:	sigmoid = 21'b111111111111111010011;
		14'b01010110000110:	sigmoid = 21'b111111111111111010011;
		14'b01010110000111:	sigmoid = 21'b111111111111111010011;
		14'b01010110001000:	sigmoid = 21'b111111111111111010011;
		14'b01010110001001:	sigmoid = 21'b111111111111111010011;
		14'b01010110001010:	sigmoid = 21'b111111111111111010011;
		14'b01010110001011:	sigmoid = 21'b111111111111111010011;
		14'b01010110001100:	sigmoid = 21'b111111111111111010100;
		14'b01010110001101:	sigmoid = 21'b111111111111111010100;
		14'b01010110001110:	sigmoid = 21'b111111111111111010100;
		14'b01010110001111:	sigmoid = 21'b111111111111111010100;
		14'b01010110010000:	sigmoid = 21'b111111111111111010100;
		14'b01010110010001:	sigmoid = 21'b111111111111111010100;
		14'b01010110010010:	sigmoid = 21'b111111111111111010100;
		14'b01010110010011:	sigmoid = 21'b111111111111111010100;
		14'b01010110010100:	sigmoid = 21'b111111111111111010100;
		14'b01010110010101:	sigmoid = 21'b111111111111111010100;
		14'b01010110010110:	sigmoid = 21'b111111111111111010100;
		14'b01010110010111:	sigmoid = 21'b111111111111111010101;
		14'b01010110011000:	sigmoid = 21'b111111111111111010101;
		14'b01010110011001:	sigmoid = 21'b111111111111111010101;
		14'b01010110011010:	sigmoid = 21'b111111111111111010101;
		14'b01010110011011:	sigmoid = 21'b111111111111111010101;
		14'b01010110011100:	sigmoid = 21'b111111111111111010101;
		14'b01010110011101:	sigmoid = 21'b111111111111111010101;
		14'b01010110011110:	sigmoid = 21'b111111111111111010101;
		14'b01010110011111:	sigmoid = 21'b111111111111111010101;
		14'b01010110100000:	sigmoid = 21'b111111111111111010101;
		14'b01010110100001:	sigmoid = 21'b111111111111111010101;
		14'b01010110100010:	sigmoid = 21'b111111111111111010101;
		14'b01010110100011:	sigmoid = 21'b111111111111111010101;
		14'b01010110100100:	sigmoid = 21'b111111111111111010110;
		14'b01010110100101:	sigmoid = 21'b111111111111111010110;
		14'b01010110100110:	sigmoid = 21'b111111111111111010110;
		14'b01010110100111:	sigmoid = 21'b111111111111111010110;
		14'b01010110101000:	sigmoid = 21'b111111111111111010110;
		14'b01010110101001:	sigmoid = 21'b111111111111111010110;
		14'b01010110101010:	sigmoid = 21'b111111111111111010110;
		14'b01010110101011:	sigmoid = 21'b111111111111111010110;
		14'b01010110101100:	sigmoid = 21'b111111111111111010110;
		14'b01010110101101:	sigmoid = 21'b111111111111111010110;
		14'b01010110101110:	sigmoid = 21'b111111111111111010110;
		14'b01010110101111:	sigmoid = 21'b111111111111111010110;
		14'b01010110110000:	sigmoid = 21'b111111111111111010111;
		14'b01010110110001:	sigmoid = 21'b111111111111111010111;
		14'b01010110110010:	sigmoid = 21'b111111111111111010111;
		14'b01010110110011:	sigmoid = 21'b111111111111111010111;
		14'b01010110110100:	sigmoid = 21'b111111111111111010111;
		14'b01010110110101:	sigmoid = 21'b111111111111111010111;
		14'b01010110110110:	sigmoid = 21'b111111111111111010111;
		14'b01010110110111:	sigmoid = 21'b111111111111111010111;
		14'b01010110111000:	sigmoid = 21'b111111111111111010111;
		14'b01010110111001:	sigmoid = 21'b111111111111111010111;
		14'b01010110111010:	sigmoid = 21'b111111111111111010111;
		14'b01010110111011:	sigmoid = 21'b111111111111111010111;
		14'b01010110111100:	sigmoid = 21'b111111111111111010111;
		14'b01010110111101:	sigmoid = 21'b111111111111111011000;
		14'b01010110111110:	sigmoid = 21'b111111111111111011000;
		14'b01010110111111:	sigmoid = 21'b111111111111111011000;
		14'b01010111000000:	sigmoid = 21'b111111111111111011000;
		14'b01010111000001:	sigmoid = 21'b111111111111111011000;
		14'b01010111000010:	sigmoid = 21'b111111111111111011000;
		14'b01010111000011:	sigmoid = 21'b111111111111111011000;
		14'b01010111000100:	sigmoid = 21'b111111111111111011000;
		14'b01010111000101:	sigmoid = 21'b111111111111111011000;
		14'b01010111000110:	sigmoid = 21'b111111111111111011000;
		14'b01010111000111:	sigmoid = 21'b111111111111111011000;
		14'b01010111001000:	sigmoid = 21'b111111111111111011000;
		14'b01010111001001:	sigmoid = 21'b111111111111111011001;
		14'b01010111001010:	sigmoid = 21'b111111111111111011001;
		14'b01010111001011:	sigmoid = 21'b111111111111111011001;
		14'b01010111001100:	sigmoid = 21'b111111111111111011001;
		14'b01010111001101:	sigmoid = 21'b111111111111111011001;
		14'b01010111001110:	sigmoid = 21'b111111111111111011001;
		14'b01010111001111:	sigmoid = 21'b111111111111111011001;
		14'b01010111010000:	sigmoid = 21'b111111111111111011001;
		14'b01010111010001:	sigmoid = 21'b111111111111111011001;
		14'b01010111010010:	sigmoid = 21'b111111111111111011001;
		14'b01010111010011:	sigmoid = 21'b111111111111111011001;
		14'b01010111010100:	sigmoid = 21'b111111111111111011001;
		14'b01010111010101:	sigmoid = 21'b111111111111111011001;
		14'b01010111010110:	sigmoid = 21'b111111111111111011001;
		14'b01010111010111:	sigmoid = 21'b111111111111111011010;
		14'b01010111011000:	sigmoid = 21'b111111111111111011010;
		14'b01010111011001:	sigmoid = 21'b111111111111111011010;
		14'b01010111011010:	sigmoid = 21'b111111111111111011010;
		14'b01010111011011:	sigmoid = 21'b111111111111111011010;
		14'b01010111011100:	sigmoid = 21'b111111111111111011010;
		14'b01010111011101:	sigmoid = 21'b111111111111111011010;
		14'b01010111011110:	sigmoid = 21'b111111111111111011010;
		14'b01010111011111:	sigmoid = 21'b111111111111111011010;
		14'b01010111100000:	sigmoid = 21'b111111111111111011010;
		14'b01010111100001:	sigmoid = 21'b111111111111111011010;
		14'b01010111100010:	sigmoid = 21'b111111111111111011010;
		14'b01010111100011:	sigmoid = 21'b111111111111111011010;
		14'b01010111100100:	sigmoid = 21'b111111111111111011011;
		14'b01010111100101:	sigmoid = 21'b111111111111111011011;
		14'b01010111100110:	sigmoid = 21'b111111111111111011011;
		14'b01010111100111:	sigmoid = 21'b111111111111111011011;
		14'b01010111101000:	sigmoid = 21'b111111111111111011011;
		14'b01010111101001:	sigmoid = 21'b111111111111111011011;
		14'b01010111101010:	sigmoid = 21'b111111111111111011011;
		14'b01010111101011:	sigmoid = 21'b111111111111111011011;
		14'b01010111101100:	sigmoid = 21'b111111111111111011011;
		14'b01010111101101:	sigmoid = 21'b111111111111111011011;
		14'b01010111101110:	sigmoid = 21'b111111111111111011011;
		14'b01010111101111:	sigmoid = 21'b111111111111111011011;
		14'b01010111110000:	sigmoid = 21'b111111111111111011011;
		14'b01010111110001:	sigmoid = 21'b111111111111111011011;
		14'b01010111110010:	sigmoid = 21'b111111111111111011100;
		14'b01010111110011:	sigmoid = 21'b111111111111111011100;
		14'b01010111110100:	sigmoid = 21'b111111111111111011100;
		14'b01010111110101:	sigmoid = 21'b111111111111111011100;
		14'b01010111110110:	sigmoid = 21'b111111111111111011100;
		14'b01010111110111:	sigmoid = 21'b111111111111111011100;
		14'b01010111111000:	sigmoid = 21'b111111111111111011100;
		14'b01010111111001:	sigmoid = 21'b111111111111111011100;
		14'b01010111111010:	sigmoid = 21'b111111111111111011100;
		14'b01010111111011:	sigmoid = 21'b111111111111111011100;
		14'b01010111111100:	sigmoid = 21'b111111111111111011100;
		14'b01010111111101:	sigmoid = 21'b111111111111111011100;
		14'b01010111111110:	sigmoid = 21'b111111111111111011100;
		14'b01010111111111:	sigmoid = 21'b111111111111111011100;
		14'b01011000000000:	sigmoid = 21'b111111111111111011100;
		14'b01011000000001:	sigmoid = 21'b111111111111111011101;
		14'b01011000000010:	sigmoid = 21'b111111111111111011101;
		14'b01011000000011:	sigmoid = 21'b111111111111111011101;
		14'b01011000000100:	sigmoid = 21'b111111111111111011101;
		14'b01011000000101:	sigmoid = 21'b111111111111111011101;
		14'b01011000000110:	sigmoid = 21'b111111111111111011101;
		14'b01011000000111:	sigmoid = 21'b111111111111111011101;
		14'b01011000001000:	sigmoid = 21'b111111111111111011101;
		14'b01011000001001:	sigmoid = 21'b111111111111111011101;
		14'b01011000001010:	sigmoid = 21'b111111111111111011101;
		14'b01011000001011:	sigmoid = 21'b111111111111111011101;
		14'b01011000001100:	sigmoid = 21'b111111111111111011101;
		14'b01011000001101:	sigmoid = 21'b111111111111111011101;
		14'b01011000001110:	sigmoid = 21'b111111111111111011101;
		14'b01011000001111:	sigmoid = 21'b111111111111111011101;
		14'b01011000010000:	sigmoid = 21'b111111111111111011110;
		14'b01011000010001:	sigmoid = 21'b111111111111111011110;
		14'b01011000010010:	sigmoid = 21'b111111111111111011110;
		14'b01011000010011:	sigmoid = 21'b111111111111111011110;
		14'b01011000010100:	sigmoid = 21'b111111111111111011110;
		14'b01011000010101:	sigmoid = 21'b111111111111111011110;
		14'b01011000010110:	sigmoid = 21'b111111111111111011110;
		14'b01011000010111:	sigmoid = 21'b111111111111111011110;
		14'b01011000011000:	sigmoid = 21'b111111111111111011110;
		14'b01011000011001:	sigmoid = 21'b111111111111111011110;
		14'b01011000011010:	sigmoid = 21'b111111111111111011110;
		14'b01011000011011:	sigmoid = 21'b111111111111111011110;
		14'b01011000011100:	sigmoid = 21'b111111111111111011110;
		14'b01011000011101:	sigmoid = 21'b111111111111111011110;
		14'b01011000011110:	sigmoid = 21'b111111111111111011110;
		14'b01011000011111:	sigmoid = 21'b111111111111111011111;
		14'b01011000100000:	sigmoid = 21'b111111111111111011111;
		14'b01011000100001:	sigmoid = 21'b111111111111111011111;
		14'b01011000100010:	sigmoid = 21'b111111111111111011111;
		14'b01011000100011:	sigmoid = 21'b111111111111111011111;
		14'b01011000100100:	sigmoid = 21'b111111111111111011111;
		14'b01011000100101:	sigmoid = 21'b111111111111111011111;
		14'b01011000100110:	sigmoid = 21'b111111111111111011111;
		14'b01011000100111:	sigmoid = 21'b111111111111111011111;
		14'b01011000101000:	sigmoid = 21'b111111111111111011111;
		14'b01011000101001:	sigmoid = 21'b111111111111111011111;
		14'b01011000101010:	sigmoid = 21'b111111111111111011111;
		14'b01011000101011:	sigmoid = 21'b111111111111111011111;
		14'b01011000101100:	sigmoid = 21'b111111111111111011111;
		14'b01011000101101:	sigmoid = 21'b111111111111111011111;
		14'b01011000101110:	sigmoid = 21'b111111111111111011111;
		14'b01011000101111:	sigmoid = 21'b111111111111111100000;
		14'b01011000110000:	sigmoid = 21'b111111111111111100000;
		14'b01011000110001:	sigmoid = 21'b111111111111111100000;
		14'b01011000110010:	sigmoid = 21'b111111111111111100000;
		14'b01011000110011:	sigmoid = 21'b111111111111111100000;
		14'b01011000110100:	sigmoid = 21'b111111111111111100000;
		14'b01011000110101:	sigmoid = 21'b111111111111111100000;
		14'b01011000110110:	sigmoid = 21'b111111111111111100000;
		14'b01011000110111:	sigmoid = 21'b111111111111111100000;
		14'b01011000111000:	sigmoid = 21'b111111111111111100000;
		14'b01011000111001:	sigmoid = 21'b111111111111111100000;
		14'b01011000111010:	sigmoid = 21'b111111111111111100000;
		14'b01011000111011:	sigmoid = 21'b111111111111111100000;
		14'b01011000111100:	sigmoid = 21'b111111111111111100000;
		14'b01011000111101:	sigmoid = 21'b111111111111111100000;
		14'b01011000111110:	sigmoid = 21'b111111111111111100000;
		14'b01011000111111:	sigmoid = 21'b111111111111111100001;
		14'b01011001000000:	sigmoid = 21'b111111111111111100001;
		14'b01011001000001:	sigmoid = 21'b111111111111111100001;
		14'b01011001000010:	sigmoid = 21'b111111111111111100001;
		14'b01011001000011:	sigmoid = 21'b111111111111111100001;
		14'b01011001000100:	sigmoid = 21'b111111111111111100001;
		14'b01011001000101:	sigmoid = 21'b111111111111111100001;
		14'b01011001000110:	sigmoid = 21'b111111111111111100001;
		14'b01011001000111:	sigmoid = 21'b111111111111111100001;
		14'b01011001001000:	sigmoid = 21'b111111111111111100001;
		14'b01011001001001:	sigmoid = 21'b111111111111111100001;
		14'b01011001001010:	sigmoid = 21'b111111111111111100001;
		14'b01011001001011:	sigmoid = 21'b111111111111111100001;
		14'b01011001001100:	sigmoid = 21'b111111111111111100001;
		14'b01011001001101:	sigmoid = 21'b111111111111111100001;
		14'b01011001001110:	sigmoid = 21'b111111111111111100001;
		14'b01011001001111:	sigmoid = 21'b111111111111111100001;
		14'b01011001010000:	sigmoid = 21'b111111111111111100010;
		14'b01011001010001:	sigmoid = 21'b111111111111111100010;
		14'b01011001010010:	sigmoid = 21'b111111111111111100010;
		14'b01011001010011:	sigmoid = 21'b111111111111111100010;
		14'b01011001010100:	sigmoid = 21'b111111111111111100010;
		14'b01011001010101:	sigmoid = 21'b111111111111111100010;
		14'b01011001010110:	sigmoid = 21'b111111111111111100010;
		14'b01011001010111:	sigmoid = 21'b111111111111111100010;
		14'b01011001011000:	sigmoid = 21'b111111111111111100010;
		14'b01011001011001:	sigmoid = 21'b111111111111111100010;
		14'b01011001011010:	sigmoid = 21'b111111111111111100010;
		14'b01011001011011:	sigmoid = 21'b111111111111111100010;
		14'b01011001011100:	sigmoid = 21'b111111111111111100010;
		14'b01011001011101:	sigmoid = 21'b111111111111111100010;
		14'b01011001011110:	sigmoid = 21'b111111111111111100010;
		14'b01011001011111:	sigmoid = 21'b111111111111111100010;
		14'b01011001100000:	sigmoid = 21'b111111111111111100010;
		14'b01011001100001:	sigmoid = 21'b111111111111111100011;
		14'b01011001100010:	sigmoid = 21'b111111111111111100011;
		14'b01011001100011:	sigmoid = 21'b111111111111111100011;
		14'b01011001100100:	sigmoid = 21'b111111111111111100011;
		14'b01011001100101:	sigmoid = 21'b111111111111111100011;
		14'b01011001100110:	sigmoid = 21'b111111111111111100011;
		14'b01011001100111:	sigmoid = 21'b111111111111111100011;
		14'b01011001101000:	sigmoid = 21'b111111111111111100011;
		14'b01011001101001:	sigmoid = 21'b111111111111111100011;
		14'b01011001101010:	sigmoid = 21'b111111111111111100011;
		14'b01011001101011:	sigmoid = 21'b111111111111111100011;
		14'b01011001101100:	sigmoid = 21'b111111111111111100011;
		14'b01011001101101:	sigmoid = 21'b111111111111111100011;
		14'b01011001101110:	sigmoid = 21'b111111111111111100011;
		14'b01011001101111:	sigmoid = 21'b111111111111111100011;
		14'b01011001110000:	sigmoid = 21'b111111111111111100011;
		14'b01011001110001:	sigmoid = 21'b111111111111111100011;
		14'b01011001110010:	sigmoid = 21'b111111111111111100011;
		14'b01011001110011:	sigmoid = 21'b111111111111111100100;
		14'b01011001110100:	sigmoid = 21'b111111111111111100100;
		14'b01011001110101:	sigmoid = 21'b111111111111111100100;
		14'b01011001110110:	sigmoid = 21'b111111111111111100100;
		14'b01011001110111:	sigmoid = 21'b111111111111111100100;
		14'b01011001111000:	sigmoid = 21'b111111111111111100100;
		14'b01011001111001:	sigmoid = 21'b111111111111111100100;
		14'b01011001111010:	sigmoid = 21'b111111111111111100100;
		14'b01011001111011:	sigmoid = 21'b111111111111111100100;
		14'b01011001111100:	sigmoid = 21'b111111111111111100100;
		14'b01011001111101:	sigmoid = 21'b111111111111111100100;
		14'b01011001111110:	sigmoid = 21'b111111111111111100100;
		14'b01011001111111:	sigmoid = 21'b111111111111111100100;
		14'b01011010000000:	sigmoid = 21'b111111111111111100100;
		14'b01011010000001:	sigmoid = 21'b111111111111111100100;
		14'b01011010000010:	sigmoid = 21'b111111111111111100100;
		14'b01011010000011:	sigmoid = 21'b111111111111111100100;
		14'b01011010000100:	sigmoid = 21'b111111111111111100100;
		14'b01011010000101:	sigmoid = 21'b111111111111111100100;
		14'b01011010000110:	sigmoid = 21'b111111111111111100101;
		14'b01011010000111:	sigmoid = 21'b111111111111111100101;
		14'b01011010001000:	sigmoid = 21'b111111111111111100101;
		14'b01011010001001:	sigmoid = 21'b111111111111111100101;
		14'b01011010001010:	sigmoid = 21'b111111111111111100101;
		14'b01011010001011:	sigmoid = 21'b111111111111111100101;
		14'b01011010001100:	sigmoid = 21'b111111111111111100101;
		14'b01011010001101:	sigmoid = 21'b111111111111111100101;
		14'b01011010001110:	sigmoid = 21'b111111111111111100101;
		14'b01011010001111:	sigmoid = 21'b111111111111111100101;
		14'b01011010010000:	sigmoid = 21'b111111111111111100101;
		14'b01011010010001:	sigmoid = 21'b111111111111111100101;
		14'b01011010010010:	sigmoid = 21'b111111111111111100101;
		14'b01011010010011:	sigmoid = 21'b111111111111111100101;
		14'b01011010010100:	sigmoid = 21'b111111111111111100101;
		14'b01011010010101:	sigmoid = 21'b111111111111111100101;
		14'b01011010010110:	sigmoid = 21'b111111111111111100101;
		14'b01011010010111:	sigmoid = 21'b111111111111111100101;
		14'b01011010011000:	sigmoid = 21'b111111111111111100101;
		14'b01011010011001:	sigmoid = 21'b111111111111111100110;
		14'b01011010011010:	sigmoid = 21'b111111111111111100110;
		14'b01011010011011:	sigmoid = 21'b111111111111111100110;
		14'b01011010011100:	sigmoid = 21'b111111111111111100110;
		14'b01011010011101:	sigmoid = 21'b111111111111111100110;
		14'b01011010011110:	sigmoid = 21'b111111111111111100110;
		14'b01011010011111:	sigmoid = 21'b111111111111111100110;
		14'b01011010100000:	sigmoid = 21'b111111111111111100110;
		14'b01011010100001:	sigmoid = 21'b111111111111111100110;
		14'b01011010100010:	sigmoid = 21'b111111111111111100110;
		14'b01011010100011:	sigmoid = 21'b111111111111111100110;
		14'b01011010100100:	sigmoid = 21'b111111111111111100110;
		14'b01011010100101:	sigmoid = 21'b111111111111111100110;
		14'b01011010100110:	sigmoid = 21'b111111111111111100110;
		14'b01011010100111:	sigmoid = 21'b111111111111111100110;
		14'b01011010101000:	sigmoid = 21'b111111111111111100110;
		14'b01011010101001:	sigmoid = 21'b111111111111111100110;
		14'b01011010101010:	sigmoid = 21'b111111111111111100110;
		14'b01011010101011:	sigmoid = 21'b111111111111111100110;
		14'b01011010101100:	sigmoid = 21'b111111111111111100110;
		14'b01011010101101:	sigmoid = 21'b111111111111111100111;
		14'b01011010101110:	sigmoid = 21'b111111111111111100111;
		14'b01011010101111:	sigmoid = 21'b111111111111111100111;
		14'b01011010110000:	sigmoid = 21'b111111111111111100111;
		14'b01011010110001:	sigmoid = 21'b111111111111111100111;
		14'b01011010110010:	sigmoid = 21'b111111111111111100111;
		14'b01011010110011:	sigmoid = 21'b111111111111111100111;
		14'b01011010110100:	sigmoid = 21'b111111111111111100111;
		14'b01011010110101:	sigmoid = 21'b111111111111111100111;
		14'b01011010110110:	sigmoid = 21'b111111111111111100111;
		14'b01011010110111:	sigmoid = 21'b111111111111111100111;
		14'b01011010111000:	sigmoid = 21'b111111111111111100111;
		14'b01011010111001:	sigmoid = 21'b111111111111111100111;
		14'b01011010111010:	sigmoid = 21'b111111111111111100111;
		14'b01011010111011:	sigmoid = 21'b111111111111111100111;
		14'b01011010111100:	sigmoid = 21'b111111111111111100111;
		14'b01011010111101:	sigmoid = 21'b111111111111111100111;
		14'b01011010111110:	sigmoid = 21'b111111111111111100111;
		14'b01011010111111:	sigmoid = 21'b111111111111111100111;
		14'b01011011000000:	sigmoid = 21'b111111111111111100111;
		14'b01011011000001:	sigmoid = 21'b111111111111111100111;
		14'b01011011000010:	sigmoid = 21'b111111111111111101000;
		14'b01011011000011:	sigmoid = 21'b111111111111111101000;
		14'b01011011000100:	sigmoid = 21'b111111111111111101000;
		14'b01011011000101:	sigmoid = 21'b111111111111111101000;
		14'b01011011000110:	sigmoid = 21'b111111111111111101000;
		14'b01011011000111:	sigmoid = 21'b111111111111111101000;
		14'b01011011001000:	sigmoid = 21'b111111111111111101000;
		14'b01011011001001:	sigmoid = 21'b111111111111111101000;
		14'b01011011001010:	sigmoid = 21'b111111111111111101000;
		14'b01011011001011:	sigmoid = 21'b111111111111111101000;
		14'b01011011001100:	sigmoid = 21'b111111111111111101000;
		14'b01011011001101:	sigmoid = 21'b111111111111111101000;
		14'b01011011001110:	sigmoid = 21'b111111111111111101000;
		14'b01011011001111:	sigmoid = 21'b111111111111111101000;
		14'b01011011010000:	sigmoid = 21'b111111111111111101000;
		14'b01011011010001:	sigmoid = 21'b111111111111111101000;
		14'b01011011010010:	sigmoid = 21'b111111111111111101000;
		14'b01011011010011:	sigmoid = 21'b111111111111111101000;
		14'b01011011010100:	sigmoid = 21'b111111111111111101000;
		14'b01011011010101:	sigmoid = 21'b111111111111111101000;
		14'b01011011010110:	sigmoid = 21'b111111111111111101000;
		14'b01011011010111:	sigmoid = 21'b111111111111111101000;
		14'b01011011011000:	sigmoid = 21'b111111111111111101001;
		14'b01011011011001:	sigmoid = 21'b111111111111111101001;
		14'b01011011011010:	sigmoid = 21'b111111111111111101001;
		14'b01011011011011:	sigmoid = 21'b111111111111111101001;
		14'b01011011011100:	sigmoid = 21'b111111111111111101001;
		14'b01011011011101:	sigmoid = 21'b111111111111111101001;
		14'b01011011011110:	sigmoid = 21'b111111111111111101001;
		14'b01011011011111:	sigmoid = 21'b111111111111111101001;
		14'b01011011100000:	sigmoid = 21'b111111111111111101001;
		14'b01011011100001:	sigmoid = 21'b111111111111111101001;
		14'b01011011100010:	sigmoid = 21'b111111111111111101001;
		14'b01011011100011:	sigmoid = 21'b111111111111111101001;
		14'b01011011100100:	sigmoid = 21'b111111111111111101001;
		14'b01011011100101:	sigmoid = 21'b111111111111111101001;
		14'b01011011100110:	sigmoid = 21'b111111111111111101001;
		14'b01011011100111:	sigmoid = 21'b111111111111111101001;
		14'b01011011101000:	sigmoid = 21'b111111111111111101001;
		14'b01011011101001:	sigmoid = 21'b111111111111111101001;
		14'b01011011101010:	sigmoid = 21'b111111111111111101001;
		14'b01011011101011:	sigmoid = 21'b111111111111111101001;
		14'b01011011101100:	sigmoid = 21'b111111111111111101001;
		14'b01011011101101:	sigmoid = 21'b111111111111111101001;
		14'b01011011101110:	sigmoid = 21'b111111111111111101001;
		14'b01011011101111:	sigmoid = 21'b111111111111111101010;
		14'b01011011110000:	sigmoid = 21'b111111111111111101010;
		14'b01011011110001:	sigmoid = 21'b111111111111111101010;
		14'b01011011110010:	sigmoid = 21'b111111111111111101010;
		14'b01011011110011:	sigmoid = 21'b111111111111111101010;
		14'b01011011110100:	sigmoid = 21'b111111111111111101010;
		14'b01011011110101:	sigmoid = 21'b111111111111111101010;
		14'b01011011110110:	sigmoid = 21'b111111111111111101010;
		14'b01011011110111:	sigmoid = 21'b111111111111111101010;
		14'b01011011111000:	sigmoid = 21'b111111111111111101010;
		14'b01011011111001:	sigmoid = 21'b111111111111111101010;
		14'b01011011111010:	sigmoid = 21'b111111111111111101010;
		14'b01011011111011:	sigmoid = 21'b111111111111111101010;
		14'b01011011111100:	sigmoid = 21'b111111111111111101010;
		14'b01011011111101:	sigmoid = 21'b111111111111111101010;
		14'b01011011111110:	sigmoid = 21'b111111111111111101010;
		14'b01011011111111:	sigmoid = 21'b111111111111111101010;
		14'b01011100000000:	sigmoid = 21'b111111111111111101010;
		14'b01011100000001:	sigmoid = 21'b111111111111111101010;
		14'b01011100000010:	sigmoid = 21'b111111111111111101010;
		14'b01011100000011:	sigmoid = 21'b111111111111111101010;
		14'b01011100000100:	sigmoid = 21'b111111111111111101010;
		14'b01011100000101:	sigmoid = 21'b111111111111111101010;
		14'b01011100000110:	sigmoid = 21'b111111111111111101011;
		14'b01011100000111:	sigmoid = 21'b111111111111111101011;
		14'b01011100001000:	sigmoid = 21'b111111111111111101011;
		14'b01011100001001:	sigmoid = 21'b111111111111111101011;
		14'b01011100001010:	sigmoid = 21'b111111111111111101011;
		14'b01011100001011:	sigmoid = 21'b111111111111111101011;
		14'b01011100001100:	sigmoid = 21'b111111111111111101011;
		14'b01011100001101:	sigmoid = 21'b111111111111111101011;
		14'b01011100001110:	sigmoid = 21'b111111111111111101011;
		14'b01011100001111:	sigmoid = 21'b111111111111111101011;
		14'b01011100010000:	sigmoid = 21'b111111111111111101011;
		14'b01011100010001:	sigmoid = 21'b111111111111111101011;
		14'b01011100010010:	sigmoid = 21'b111111111111111101011;
		14'b01011100010011:	sigmoid = 21'b111111111111111101011;
		14'b01011100010100:	sigmoid = 21'b111111111111111101011;
		14'b01011100010101:	sigmoid = 21'b111111111111111101011;
		14'b01011100010110:	sigmoid = 21'b111111111111111101011;
		14'b01011100010111:	sigmoid = 21'b111111111111111101011;
		14'b01011100011000:	sigmoid = 21'b111111111111111101011;
		14'b01011100011001:	sigmoid = 21'b111111111111111101011;
		14'b01011100011010:	sigmoid = 21'b111111111111111101011;
		14'b01011100011011:	sigmoid = 21'b111111111111111101011;
		14'b01011100011100:	sigmoid = 21'b111111111111111101011;
		14'b01011100011101:	sigmoid = 21'b111111111111111101011;
		14'b01011100011110:	sigmoid = 21'b111111111111111101011;
		14'b01011100011111:	sigmoid = 21'b111111111111111101100;
		14'b01011100100000:	sigmoid = 21'b111111111111111101100;
		14'b01011100100001:	sigmoid = 21'b111111111111111101100;
		14'b01011100100010:	sigmoid = 21'b111111111111111101100;
		14'b01011100100011:	sigmoid = 21'b111111111111111101100;
		14'b01011100100100:	sigmoid = 21'b111111111111111101100;
		14'b01011100100101:	sigmoid = 21'b111111111111111101100;
		14'b01011100100110:	sigmoid = 21'b111111111111111101100;
		14'b01011100100111:	sigmoid = 21'b111111111111111101100;
		14'b01011100101000:	sigmoid = 21'b111111111111111101100;
		14'b01011100101001:	sigmoid = 21'b111111111111111101100;
		14'b01011100101010:	sigmoid = 21'b111111111111111101100;
		14'b01011100101011:	sigmoid = 21'b111111111111111101100;
		14'b01011100101100:	sigmoid = 21'b111111111111111101100;
		14'b01011100101101:	sigmoid = 21'b111111111111111101100;
		14'b01011100101110:	sigmoid = 21'b111111111111111101100;
		14'b01011100101111:	sigmoid = 21'b111111111111111101100;
		14'b01011100110000:	sigmoid = 21'b111111111111111101100;
		14'b01011100110001:	sigmoid = 21'b111111111111111101100;
		14'b01011100110010:	sigmoid = 21'b111111111111111101100;
		14'b01011100110011:	sigmoid = 21'b111111111111111101100;
		14'b01011100110100:	sigmoid = 21'b111111111111111101100;
		14'b01011100110101:	sigmoid = 21'b111111111111111101100;
		14'b01011100110110:	sigmoid = 21'b111111111111111101100;
		14'b01011100110111:	sigmoid = 21'b111111111111111101100;
		14'b01011100111000:	sigmoid = 21'b111111111111111101100;
		14'b01011100111001:	sigmoid = 21'b111111111111111101100;
		14'b01011100111010:	sigmoid = 21'b111111111111111101101;
		14'b01011100111011:	sigmoid = 21'b111111111111111101101;
		14'b01011100111100:	sigmoid = 21'b111111111111111101101;
		14'b01011100111101:	sigmoid = 21'b111111111111111101101;
		14'b01011100111110:	sigmoid = 21'b111111111111111101101;
		14'b01011100111111:	sigmoid = 21'b111111111111111101101;
		14'b01011101000000:	sigmoid = 21'b111111111111111101101;
		14'b01011101000001:	sigmoid = 21'b111111111111111101101;
		14'b01011101000010:	sigmoid = 21'b111111111111111101101;
		14'b01011101000011:	sigmoid = 21'b111111111111111101101;
		14'b01011101000100:	sigmoid = 21'b111111111111111101101;
		14'b01011101000101:	sigmoid = 21'b111111111111111101101;
		14'b01011101000110:	sigmoid = 21'b111111111111111101101;
		14'b01011101000111:	sigmoid = 21'b111111111111111101101;
		14'b01011101001000:	sigmoid = 21'b111111111111111101101;
		14'b01011101001001:	sigmoid = 21'b111111111111111101101;
		14'b01011101001010:	sigmoid = 21'b111111111111111101101;
		14'b01011101001011:	sigmoid = 21'b111111111111111101101;
		14'b01011101001100:	sigmoid = 21'b111111111111111101101;
		14'b01011101001101:	sigmoid = 21'b111111111111111101101;
		14'b01011101001110:	sigmoid = 21'b111111111111111101101;
		14'b01011101001111:	sigmoid = 21'b111111111111111101101;
		14'b01011101010000:	sigmoid = 21'b111111111111111101101;
		14'b01011101010001:	sigmoid = 21'b111111111111111101101;
		14'b01011101010010:	sigmoid = 21'b111111111111111101101;
		14'b01011101010011:	sigmoid = 21'b111111111111111101101;
		14'b01011101010100:	sigmoid = 21'b111111111111111101101;
		14'b01011101010101:	sigmoid = 21'b111111111111111101110;
		14'b01011101010110:	sigmoid = 21'b111111111111111101110;
		14'b01011101010111:	sigmoid = 21'b111111111111111101110;
		14'b01011101011000:	sigmoid = 21'b111111111111111101110;
		14'b01011101011001:	sigmoid = 21'b111111111111111101110;
		14'b01011101011010:	sigmoid = 21'b111111111111111101110;
		14'b01011101011011:	sigmoid = 21'b111111111111111101110;
		14'b01011101011100:	sigmoid = 21'b111111111111111101110;
		14'b01011101011101:	sigmoid = 21'b111111111111111101110;
		14'b01011101011110:	sigmoid = 21'b111111111111111101110;
		14'b01011101011111:	sigmoid = 21'b111111111111111101110;
		14'b01011101100000:	sigmoid = 21'b111111111111111101110;
		14'b01011101100001:	sigmoid = 21'b111111111111111101110;
		14'b01011101100010:	sigmoid = 21'b111111111111111101110;
		14'b01011101100011:	sigmoid = 21'b111111111111111101110;
		14'b01011101100100:	sigmoid = 21'b111111111111111101110;
		14'b01011101100101:	sigmoid = 21'b111111111111111101110;
		14'b01011101100110:	sigmoid = 21'b111111111111111101110;
		14'b01011101100111:	sigmoid = 21'b111111111111111101110;
		14'b01011101101000:	sigmoid = 21'b111111111111111101110;
		14'b01011101101001:	sigmoid = 21'b111111111111111101110;
		14'b01011101101010:	sigmoid = 21'b111111111111111101110;
		14'b01011101101011:	sigmoid = 21'b111111111111111101110;
		14'b01011101101100:	sigmoid = 21'b111111111111111101110;
		14'b01011101101101:	sigmoid = 21'b111111111111111101110;
		14'b01011101101110:	sigmoid = 21'b111111111111111101110;
		14'b01011101101111:	sigmoid = 21'b111111111111111101110;
		14'b01011101110000:	sigmoid = 21'b111111111111111101110;
		14'b01011101110001:	sigmoid = 21'b111111111111111101110;
		14'b01011101110010:	sigmoid = 21'b111111111111111101110;
		14'b01011101110011:	sigmoid = 21'b111111111111111101111;
		14'b01011101110100:	sigmoid = 21'b111111111111111101111;
		14'b01011101110101:	sigmoid = 21'b111111111111111101111;
		14'b01011101110110:	sigmoid = 21'b111111111111111101111;
		14'b01011101110111:	sigmoid = 21'b111111111111111101111;
		14'b01011101111000:	sigmoid = 21'b111111111111111101111;
		14'b01011101111001:	sigmoid = 21'b111111111111111101111;
		14'b01011101111010:	sigmoid = 21'b111111111111111101111;
		14'b01011101111011:	sigmoid = 21'b111111111111111101111;
		14'b01011101111100:	sigmoid = 21'b111111111111111101111;
		14'b01011101111101:	sigmoid = 21'b111111111111111101111;
		14'b01011101111110:	sigmoid = 21'b111111111111111101111;
		14'b01011101111111:	sigmoid = 21'b111111111111111101111;
		14'b01011110000000:	sigmoid = 21'b111111111111111101111;
		14'b01011110000001:	sigmoid = 21'b111111111111111101111;
		14'b01011110000010:	sigmoid = 21'b111111111111111101111;
		14'b01011110000011:	sigmoid = 21'b111111111111111101111;
		14'b01011110000100:	sigmoid = 21'b111111111111111101111;
		14'b01011110000101:	sigmoid = 21'b111111111111111101111;
		14'b01011110000110:	sigmoid = 21'b111111111111111101111;
		14'b01011110000111:	sigmoid = 21'b111111111111111101111;
		14'b01011110001000:	sigmoid = 21'b111111111111111101111;
		14'b01011110001001:	sigmoid = 21'b111111111111111101111;
		14'b01011110001010:	sigmoid = 21'b111111111111111101111;
		14'b01011110001011:	sigmoid = 21'b111111111111111101111;
		14'b01011110001100:	sigmoid = 21'b111111111111111101111;
		14'b01011110001101:	sigmoid = 21'b111111111111111101111;
		14'b01011110001110:	sigmoid = 21'b111111111111111101111;
		14'b01011110001111:	sigmoid = 21'b111111111111111101111;
		14'b01011110010000:	sigmoid = 21'b111111111111111101111;
		14'b01011110010001:	sigmoid = 21'b111111111111111101111;
		14'b01011110010010:	sigmoid = 21'b111111111111111110000;
		14'b01011110010011:	sigmoid = 21'b111111111111111110000;
		14'b01011110010100:	sigmoid = 21'b111111111111111110000;
		14'b01011110010101:	sigmoid = 21'b111111111111111110000;
		14'b01011110010110:	sigmoid = 21'b111111111111111110000;
		14'b01011110010111:	sigmoid = 21'b111111111111111110000;
		14'b01011110011000:	sigmoid = 21'b111111111111111110000;
		14'b01011110011001:	sigmoid = 21'b111111111111111110000;
		14'b01011110011010:	sigmoid = 21'b111111111111111110000;
		14'b01011110011011:	sigmoid = 21'b111111111111111110000;
		14'b01011110011100:	sigmoid = 21'b111111111111111110000;
		14'b01011110011101:	sigmoid = 21'b111111111111111110000;
		14'b01011110011110:	sigmoid = 21'b111111111111111110000;
		14'b01011110011111:	sigmoid = 21'b111111111111111110000;
		14'b01011110100000:	sigmoid = 21'b111111111111111110000;
		14'b01011110100001:	sigmoid = 21'b111111111111111110000;
		14'b01011110100010:	sigmoid = 21'b111111111111111110000;
		14'b01011110100011:	sigmoid = 21'b111111111111111110000;
		14'b01011110100100:	sigmoid = 21'b111111111111111110000;
		14'b01011110100101:	sigmoid = 21'b111111111111111110000;
		14'b01011110100110:	sigmoid = 21'b111111111111111110000;
		14'b01011110100111:	sigmoid = 21'b111111111111111110000;
		14'b01011110101000:	sigmoid = 21'b111111111111111110000;
		14'b01011110101001:	sigmoid = 21'b111111111111111110000;
		14'b01011110101010:	sigmoid = 21'b111111111111111110000;
		14'b01011110101011:	sigmoid = 21'b111111111111111110000;
		14'b01011110101100:	sigmoid = 21'b111111111111111110000;
		14'b01011110101101:	sigmoid = 21'b111111111111111110000;
		14'b01011110101110:	sigmoid = 21'b111111111111111110000;
		14'b01011110101111:	sigmoid = 21'b111111111111111110000;
		14'b01011110110000:	sigmoid = 21'b111111111111111110000;
		14'b01011110110001:	sigmoid = 21'b111111111111111110000;
		14'b01011110110010:	sigmoid = 21'b111111111111111110000;
		14'b01011110110011:	sigmoid = 21'b111111111111111110001;
		14'b01011110110100:	sigmoid = 21'b111111111111111110001;
		14'b01011110110101:	sigmoid = 21'b111111111111111110001;
		14'b01011110110110:	sigmoid = 21'b111111111111111110001;
		14'b01011110110111:	sigmoid = 21'b111111111111111110001;
		14'b01011110111000:	sigmoid = 21'b111111111111111110001;
		14'b01011110111001:	sigmoid = 21'b111111111111111110001;
		14'b01011110111010:	sigmoid = 21'b111111111111111110001;
		14'b01011110111011:	sigmoid = 21'b111111111111111110001;
		14'b01011110111100:	sigmoid = 21'b111111111111111110001;
		14'b01011110111101:	sigmoid = 21'b111111111111111110001;
		14'b01011110111110:	sigmoid = 21'b111111111111111110001;
		14'b01011110111111:	sigmoid = 21'b111111111111111110001;
		14'b01011111000000:	sigmoid = 21'b111111111111111110001;
		14'b01011111000001:	sigmoid = 21'b111111111111111110001;
		14'b01011111000010:	sigmoid = 21'b111111111111111110001;
		14'b01011111000011:	sigmoid = 21'b111111111111111110001;
		14'b01011111000100:	sigmoid = 21'b111111111111111110001;
		14'b01011111000101:	sigmoid = 21'b111111111111111110001;
		14'b01011111000110:	sigmoid = 21'b111111111111111110001;
		14'b01011111000111:	sigmoid = 21'b111111111111111110001;
		14'b01011111001000:	sigmoid = 21'b111111111111111110001;
		14'b01011111001001:	sigmoid = 21'b111111111111111110001;
		14'b01011111001010:	sigmoid = 21'b111111111111111110001;
		14'b01011111001011:	sigmoid = 21'b111111111111111110001;
		14'b01011111001100:	sigmoid = 21'b111111111111111110001;
		14'b01011111001101:	sigmoid = 21'b111111111111111110001;
		14'b01011111001110:	sigmoid = 21'b111111111111111110001;
		14'b01011111001111:	sigmoid = 21'b111111111111111110001;
		14'b01011111010000:	sigmoid = 21'b111111111111111110001;
		14'b01011111010001:	sigmoid = 21'b111111111111111110001;
		14'b01011111010010:	sigmoid = 21'b111111111111111110001;
		14'b01011111010011:	sigmoid = 21'b111111111111111110001;
		14'b01011111010100:	sigmoid = 21'b111111111111111110001;
		14'b01011111010101:	sigmoid = 21'b111111111111111110001;
		14'b01011111010110:	sigmoid = 21'b111111111111111110010;
		14'b01011111010111:	sigmoid = 21'b111111111111111110010;
		14'b01011111011000:	sigmoid = 21'b111111111111111110010;
		14'b01011111011001:	sigmoid = 21'b111111111111111110010;
		14'b01011111011010:	sigmoid = 21'b111111111111111110010;
		14'b01011111011011:	sigmoid = 21'b111111111111111110010;
		14'b01011111011100:	sigmoid = 21'b111111111111111110010;
		14'b01011111011101:	sigmoid = 21'b111111111111111110010;
		14'b01011111011110:	sigmoid = 21'b111111111111111110010;
		14'b01011111011111:	sigmoid = 21'b111111111111111110010;
		14'b01011111100000:	sigmoid = 21'b111111111111111110010;
		14'b01011111100001:	sigmoid = 21'b111111111111111110010;
		14'b01011111100010:	sigmoid = 21'b111111111111111110010;
		14'b01011111100011:	sigmoid = 21'b111111111111111110010;
		14'b01011111100100:	sigmoid = 21'b111111111111111110010;
		14'b01011111100101:	sigmoid = 21'b111111111111111110010;
		14'b01011111100110:	sigmoid = 21'b111111111111111110010;
		14'b01011111100111:	sigmoid = 21'b111111111111111110010;
		14'b01011111101000:	sigmoid = 21'b111111111111111110010;
		14'b01011111101001:	sigmoid = 21'b111111111111111110010;
		14'b01011111101010:	sigmoid = 21'b111111111111111110010;
		14'b01011111101011:	sigmoid = 21'b111111111111111110010;
		14'b01011111101100:	sigmoid = 21'b111111111111111110010;
		14'b01011111101101:	sigmoid = 21'b111111111111111110010;
		14'b01011111101110:	sigmoid = 21'b111111111111111110010;
		14'b01011111101111:	sigmoid = 21'b111111111111111110010;
		14'b01011111110000:	sigmoid = 21'b111111111111111110010;
		14'b01011111110001:	sigmoid = 21'b111111111111111110010;
		14'b01011111110010:	sigmoid = 21'b111111111111111110010;
		14'b01011111110011:	sigmoid = 21'b111111111111111110010;
		14'b01011111110100:	sigmoid = 21'b111111111111111110010;
		14'b01011111110101:	sigmoid = 21'b111111111111111110010;
		14'b01011111110110:	sigmoid = 21'b111111111111111110010;
		14'b01011111110111:	sigmoid = 21'b111111111111111110010;
		14'b01011111111000:	sigmoid = 21'b111111111111111110010;
		14'b01011111111001:	sigmoid = 21'b111111111111111110010;
		14'b01011111111010:	sigmoid = 21'b111111111111111110010;
		14'b01011111111011:	sigmoid = 21'b111111111111111110010;
		14'b01011111111100:	sigmoid = 21'b111111111111111110011;
		14'b01011111111101:	sigmoid = 21'b111111111111111110011;
		14'b01011111111110:	sigmoid = 21'b111111111111111110011;
		14'b01011111111111:	sigmoid = 21'b111111111111111110011;
		14'b01100000000000:	sigmoid = 21'b111111111111111110011;
		14'b01100000000001:	sigmoid = 21'b111111111111111110011;
		14'b01100000000010:	sigmoid = 21'b111111111111111110011;
		14'b01100000000011:	sigmoid = 21'b111111111111111110011;
		14'b01100000000100:	sigmoid = 21'b111111111111111110011;
		14'b01100000000101:	sigmoid = 21'b111111111111111110011;
		14'b01100000000110:	sigmoid = 21'b111111111111111110011;
		14'b01100000000111:	sigmoid = 21'b111111111111111110011;
		14'b01100000001000:	sigmoid = 21'b111111111111111110011;
		14'b01100000001001:	sigmoid = 21'b111111111111111110011;
		14'b01100000001010:	sigmoid = 21'b111111111111111110011;
		14'b01100000001011:	sigmoid = 21'b111111111111111110011;
		14'b01100000001100:	sigmoid = 21'b111111111111111110011;
		14'b01100000001101:	sigmoid = 21'b111111111111111110011;
		14'b01100000001110:	sigmoid = 21'b111111111111111110011;
		14'b01100000001111:	sigmoid = 21'b111111111111111110011;
		14'b01100000010000:	sigmoid = 21'b111111111111111110011;
		14'b01100000010001:	sigmoid = 21'b111111111111111110011;
		14'b01100000010010:	sigmoid = 21'b111111111111111110011;
		14'b01100000010011:	sigmoid = 21'b111111111111111110011;
		14'b01100000010100:	sigmoid = 21'b111111111111111110011;
		14'b01100000010101:	sigmoid = 21'b111111111111111110011;
		14'b01100000010110:	sigmoid = 21'b111111111111111110011;
		14'b01100000010111:	sigmoid = 21'b111111111111111110011;
		14'b01100000011000:	sigmoid = 21'b111111111111111110011;
		14'b01100000011001:	sigmoid = 21'b111111111111111110011;
		14'b01100000011010:	sigmoid = 21'b111111111111111110011;
		14'b01100000011011:	sigmoid = 21'b111111111111111110011;
		14'b01100000011100:	sigmoid = 21'b111111111111111110011;
		14'b01100000011101:	sigmoid = 21'b111111111111111110011;
		14'b01100000011110:	sigmoid = 21'b111111111111111110011;
		14'b01100000011111:	sigmoid = 21'b111111111111111110011;
		14'b01100000100000:	sigmoid = 21'b111111111111111110011;
		14'b01100000100001:	sigmoid = 21'b111111111111111110011;
		14'b01100000100010:	sigmoid = 21'b111111111111111110011;
		14'b01100000100011:	sigmoid = 21'b111111111111111110011;
		14'b01100000100100:	sigmoid = 21'b111111111111111110011;
		14'b01100000100101:	sigmoid = 21'b111111111111111110100;
		14'b01100000100110:	sigmoid = 21'b111111111111111110100;
		14'b01100000100111:	sigmoid = 21'b111111111111111110100;
		14'b01100000101000:	sigmoid = 21'b111111111111111110100;
		14'b01100000101001:	sigmoid = 21'b111111111111111110100;
		14'b01100000101010:	sigmoid = 21'b111111111111111110100;
		14'b01100000101011:	sigmoid = 21'b111111111111111110100;
		14'b01100000101100:	sigmoid = 21'b111111111111111110100;
		14'b01100000101101:	sigmoid = 21'b111111111111111110100;
		14'b01100000101110:	sigmoid = 21'b111111111111111110100;
		14'b01100000101111:	sigmoid = 21'b111111111111111110100;
		14'b01100000110000:	sigmoid = 21'b111111111111111110100;
		14'b01100000110001:	sigmoid = 21'b111111111111111110100;
		14'b01100000110010:	sigmoid = 21'b111111111111111110100;
		14'b01100000110011:	sigmoid = 21'b111111111111111110100;
		14'b01100000110100:	sigmoid = 21'b111111111111111110100;
		14'b01100000110101:	sigmoid = 21'b111111111111111110100;
		14'b01100000110110:	sigmoid = 21'b111111111111111110100;
		14'b01100000110111:	sigmoid = 21'b111111111111111110100;
		14'b01100000111000:	sigmoid = 21'b111111111111111110100;
		14'b01100000111001:	sigmoid = 21'b111111111111111110100;
		14'b01100000111010:	sigmoid = 21'b111111111111111110100;
		14'b01100000111011:	sigmoid = 21'b111111111111111110100;
		14'b01100000111100:	sigmoid = 21'b111111111111111110100;
		14'b01100000111101:	sigmoid = 21'b111111111111111110100;
		14'b01100000111110:	sigmoid = 21'b111111111111111110100;
		14'b01100000111111:	sigmoid = 21'b111111111111111110100;
		14'b01100001000000:	sigmoid = 21'b111111111111111110100;
		14'b01100001000001:	sigmoid = 21'b111111111111111110100;
		14'b01100001000010:	sigmoid = 21'b111111111111111110100;
		14'b01100001000011:	sigmoid = 21'b111111111111111110100;
		14'b01100001000100:	sigmoid = 21'b111111111111111110100;
		14'b01100001000101:	sigmoid = 21'b111111111111111110100;
		14'b01100001000110:	sigmoid = 21'b111111111111111110100;
		14'b01100001000111:	sigmoid = 21'b111111111111111110100;
		14'b01100001001000:	sigmoid = 21'b111111111111111110100;
		14'b01100001001001:	sigmoid = 21'b111111111111111110100;
		14'b01100001001010:	sigmoid = 21'b111111111111111110100;
		14'b01100001001011:	sigmoid = 21'b111111111111111110100;
		14'b01100001001100:	sigmoid = 21'b111111111111111110100;
		14'b01100001001101:	sigmoid = 21'b111111111111111110100;
		14'b01100001001110:	sigmoid = 21'b111111111111111110100;
		14'b01100001001111:	sigmoid = 21'b111111111111111110100;
		14'b01100001010000:	sigmoid = 21'b111111111111111110100;
		14'b01100001010001:	sigmoid = 21'b111111111111111110101;
		14'b01100001010010:	sigmoid = 21'b111111111111111110101;
		14'b01100001010011:	sigmoid = 21'b111111111111111110101;
		14'b01100001010100:	sigmoid = 21'b111111111111111110101;
		14'b01100001010101:	sigmoid = 21'b111111111111111110101;
		14'b01100001010110:	sigmoid = 21'b111111111111111110101;
		14'b01100001010111:	sigmoid = 21'b111111111111111110101;
		14'b01100001011000:	sigmoid = 21'b111111111111111110101;
		14'b01100001011001:	sigmoid = 21'b111111111111111110101;
		14'b01100001011010:	sigmoid = 21'b111111111111111110101;
		14'b01100001011011:	sigmoid = 21'b111111111111111110101;
		14'b01100001011100:	sigmoid = 21'b111111111111111110101;
		14'b01100001011101:	sigmoid = 21'b111111111111111110101;
		14'b01100001011110:	sigmoid = 21'b111111111111111110101;
		14'b01100001011111:	sigmoid = 21'b111111111111111110101;
		14'b01100001100000:	sigmoid = 21'b111111111111111110101;
		14'b01100001100001:	sigmoid = 21'b111111111111111110101;
		14'b01100001100010:	sigmoid = 21'b111111111111111110101;
		14'b01100001100011:	sigmoid = 21'b111111111111111110101;
		14'b01100001100100:	sigmoid = 21'b111111111111111110101;
		14'b01100001100101:	sigmoid = 21'b111111111111111110101;
		14'b01100001100110:	sigmoid = 21'b111111111111111110101;
		14'b01100001100111:	sigmoid = 21'b111111111111111110101;
		14'b01100001101000:	sigmoid = 21'b111111111111111110101;
		14'b01100001101001:	sigmoid = 21'b111111111111111110101;
		14'b01100001101010:	sigmoid = 21'b111111111111111110101;
		14'b01100001101011:	sigmoid = 21'b111111111111111110101;
		14'b01100001101100:	sigmoid = 21'b111111111111111110101;
		14'b01100001101101:	sigmoid = 21'b111111111111111110101;
		14'b01100001101110:	sigmoid = 21'b111111111111111110101;
		14'b01100001101111:	sigmoid = 21'b111111111111111110101;
		14'b01100001110000:	sigmoid = 21'b111111111111111110101;
		14'b01100001110001:	sigmoid = 21'b111111111111111110101;
		14'b01100001110010:	sigmoid = 21'b111111111111111110101;
		14'b01100001110011:	sigmoid = 21'b111111111111111110101;
		14'b01100001110100:	sigmoid = 21'b111111111111111110101;
		14'b01100001110101:	sigmoid = 21'b111111111111111110101;
		14'b01100001110110:	sigmoid = 21'b111111111111111110101;
		14'b01100001110111:	sigmoid = 21'b111111111111111110101;
		14'b01100001111000:	sigmoid = 21'b111111111111111110101;
		14'b01100001111001:	sigmoid = 21'b111111111111111110101;
		14'b01100001111010:	sigmoid = 21'b111111111111111110101;
		14'b01100001111011:	sigmoid = 21'b111111111111111110101;
		14'b01100001111100:	sigmoid = 21'b111111111111111110101;
		14'b01100001111101:	sigmoid = 21'b111111111111111110101;
		14'b01100001111110:	sigmoid = 21'b111111111111111110101;
		14'b01100001111111:	sigmoid = 21'b111111111111111110101;
		14'b01100010000000:	sigmoid = 21'b111111111111111110101;
		14'b01100010000001:	sigmoid = 21'b111111111111111110101;
		14'b01100010000010:	sigmoid = 21'b111111111111111110110;
		14'b01100010000011:	sigmoid = 21'b111111111111111110110;
		14'b01100010000100:	sigmoid = 21'b111111111111111110110;
		14'b01100010000101:	sigmoid = 21'b111111111111111110110;
		14'b01100010000110:	sigmoid = 21'b111111111111111110110;
		14'b01100010000111:	sigmoid = 21'b111111111111111110110;
		14'b01100010001000:	sigmoid = 21'b111111111111111110110;
		14'b01100010001001:	sigmoid = 21'b111111111111111110110;
		14'b01100010001010:	sigmoid = 21'b111111111111111110110;
		14'b01100010001011:	sigmoid = 21'b111111111111111110110;
		14'b01100010001100:	sigmoid = 21'b111111111111111110110;
		14'b01100010001101:	sigmoid = 21'b111111111111111110110;
		14'b01100010001110:	sigmoid = 21'b111111111111111110110;
		14'b01100010001111:	sigmoid = 21'b111111111111111110110;
		14'b01100010010000:	sigmoid = 21'b111111111111111110110;
		14'b01100010010001:	sigmoid = 21'b111111111111111110110;
		14'b01100010010010:	sigmoid = 21'b111111111111111110110;
		14'b01100010010011:	sigmoid = 21'b111111111111111110110;
		14'b01100010010100:	sigmoid = 21'b111111111111111110110;
		14'b01100010010101:	sigmoid = 21'b111111111111111110110;
		14'b01100010010110:	sigmoid = 21'b111111111111111110110;
		14'b01100010010111:	sigmoid = 21'b111111111111111110110;
		14'b01100010011000:	sigmoid = 21'b111111111111111110110;
		14'b01100010011001:	sigmoid = 21'b111111111111111110110;
		14'b01100010011010:	sigmoid = 21'b111111111111111110110;
		14'b01100010011011:	sigmoid = 21'b111111111111111110110;
		14'b01100010011100:	sigmoid = 21'b111111111111111110110;
		14'b01100010011101:	sigmoid = 21'b111111111111111110110;
		14'b01100010011110:	sigmoid = 21'b111111111111111110110;
		14'b01100010011111:	sigmoid = 21'b111111111111111110110;
		14'b01100010100000:	sigmoid = 21'b111111111111111110110;
		14'b01100010100001:	sigmoid = 21'b111111111111111110110;
		14'b01100010100010:	sigmoid = 21'b111111111111111110110;
		14'b01100010100011:	sigmoid = 21'b111111111111111110110;
		14'b01100010100100:	sigmoid = 21'b111111111111111110110;
		14'b01100010100101:	sigmoid = 21'b111111111111111110110;
		14'b01100010100110:	sigmoid = 21'b111111111111111110110;
		14'b01100010100111:	sigmoid = 21'b111111111111111110110;
		14'b01100010101000:	sigmoid = 21'b111111111111111110110;
		14'b01100010101001:	sigmoid = 21'b111111111111111110110;
		14'b01100010101010:	sigmoid = 21'b111111111111111110110;
		14'b01100010101011:	sigmoid = 21'b111111111111111110110;
		14'b01100010101100:	sigmoid = 21'b111111111111111110110;
		14'b01100010101101:	sigmoid = 21'b111111111111111110110;
		14'b01100010101110:	sigmoid = 21'b111111111111111110110;
		14'b01100010101111:	sigmoid = 21'b111111111111111110110;
		14'b01100010110000:	sigmoid = 21'b111111111111111110110;
		14'b01100010110001:	sigmoid = 21'b111111111111111110110;
		14'b01100010110010:	sigmoid = 21'b111111111111111110110;
		14'b01100010110011:	sigmoid = 21'b111111111111111110110;
		14'b01100010110100:	sigmoid = 21'b111111111111111110110;
		14'b01100010110101:	sigmoid = 21'b111111111111111110110;
		14'b01100010110110:	sigmoid = 21'b111111111111111110110;
		14'b01100010110111:	sigmoid = 21'b111111111111111110110;
		14'b01100010111000:	sigmoid = 21'b111111111111111110111;
		14'b01100010111001:	sigmoid = 21'b111111111111111110111;
		14'b01100010111010:	sigmoid = 21'b111111111111111110111;
		14'b01100010111011:	sigmoid = 21'b111111111111111110111;
		14'b01100010111100:	sigmoid = 21'b111111111111111110111;
		14'b01100010111101:	sigmoid = 21'b111111111111111110111;
		14'b01100010111110:	sigmoid = 21'b111111111111111110111;
		14'b01100010111111:	sigmoid = 21'b111111111111111110111;
		14'b01100011000000:	sigmoid = 21'b111111111111111110111;
		14'b01100011000001:	sigmoid = 21'b111111111111111110111;
		14'b01100011000010:	sigmoid = 21'b111111111111111110111;
		14'b01100011000011:	sigmoid = 21'b111111111111111110111;
		14'b01100011000100:	sigmoid = 21'b111111111111111110111;
		14'b01100011000101:	sigmoid = 21'b111111111111111110111;
		14'b01100011000110:	sigmoid = 21'b111111111111111110111;
		14'b01100011000111:	sigmoid = 21'b111111111111111110111;
		14'b01100011001000:	sigmoid = 21'b111111111111111110111;
		14'b01100011001001:	sigmoid = 21'b111111111111111110111;
		14'b01100011001010:	sigmoid = 21'b111111111111111110111;
		14'b01100011001011:	sigmoid = 21'b111111111111111110111;
		14'b01100011001100:	sigmoid = 21'b111111111111111110111;
		14'b01100011001101:	sigmoid = 21'b111111111111111110111;
		14'b01100011001110:	sigmoid = 21'b111111111111111110111;
		14'b01100011001111:	sigmoid = 21'b111111111111111110111;
		14'b01100011010000:	sigmoid = 21'b111111111111111110111;
		14'b01100011010001:	sigmoid = 21'b111111111111111110111;
		14'b01100011010010:	sigmoid = 21'b111111111111111110111;
		14'b01100011010011:	sigmoid = 21'b111111111111111110111;
		14'b01100011010100:	sigmoid = 21'b111111111111111110111;
		14'b01100011010101:	sigmoid = 21'b111111111111111110111;
		14'b01100011010110:	sigmoid = 21'b111111111111111110111;
		14'b01100011010111:	sigmoid = 21'b111111111111111110111;
		14'b01100011011000:	sigmoid = 21'b111111111111111110111;
		14'b01100011011001:	sigmoid = 21'b111111111111111110111;
		14'b01100011011010:	sigmoid = 21'b111111111111111110111;
		14'b01100011011011:	sigmoid = 21'b111111111111111110111;
		14'b01100011011100:	sigmoid = 21'b111111111111111110111;
		14'b01100011011101:	sigmoid = 21'b111111111111111110111;
		14'b01100011011110:	sigmoid = 21'b111111111111111110111;
		14'b01100011011111:	sigmoid = 21'b111111111111111110111;
		14'b01100011100000:	sigmoid = 21'b111111111111111110111;
		14'b01100011100001:	sigmoid = 21'b111111111111111110111;
		14'b01100011100010:	sigmoid = 21'b111111111111111110111;
		14'b01100011100011:	sigmoid = 21'b111111111111111110111;
		14'b01100011100100:	sigmoid = 21'b111111111111111110111;
		14'b01100011100101:	sigmoid = 21'b111111111111111110111;
		14'b01100011100110:	sigmoid = 21'b111111111111111110111;
		14'b01100011100111:	sigmoid = 21'b111111111111111110111;
		14'b01100011101000:	sigmoid = 21'b111111111111111110111;
		14'b01100011101001:	sigmoid = 21'b111111111111111110111;
		14'b01100011101010:	sigmoid = 21'b111111111111111110111;
		14'b01100011101011:	sigmoid = 21'b111111111111111110111;
		14'b01100011101100:	sigmoid = 21'b111111111111111110111;
		14'b01100011101101:	sigmoid = 21'b111111111111111110111;
		14'b01100011101110:	sigmoid = 21'b111111111111111110111;
		14'b01100011101111:	sigmoid = 21'b111111111111111110111;
		14'b01100011110000:	sigmoid = 21'b111111111111111110111;
		14'b01100011110001:	sigmoid = 21'b111111111111111110111;
		14'b01100011110010:	sigmoid = 21'b111111111111111110111;
		14'b01100011110011:	sigmoid = 21'b111111111111111110111;
		14'b01100011110100:	sigmoid = 21'b111111111111111110111;
		14'b01100011110101:	sigmoid = 21'b111111111111111111000;
		14'b01100011110110:	sigmoid = 21'b111111111111111111000;
		14'b01100011110111:	sigmoid = 21'b111111111111111111000;
		14'b01100011111000:	sigmoid = 21'b111111111111111111000;
		14'b01100011111001:	sigmoid = 21'b111111111111111111000;
		14'b01100011111010:	sigmoid = 21'b111111111111111111000;
		14'b01100011111011:	sigmoid = 21'b111111111111111111000;
		14'b01100011111100:	sigmoid = 21'b111111111111111111000;
		14'b01100011111101:	sigmoid = 21'b111111111111111111000;
		14'b01100011111110:	sigmoid = 21'b111111111111111111000;
		14'b01100011111111:	sigmoid = 21'b111111111111111111000;
		14'b01100100000000:	sigmoid = 21'b111111111111111111000;
		14'b01100100000001:	sigmoid = 21'b111111111111111111000;
		14'b01100100000010:	sigmoid = 21'b111111111111111111000;
		14'b01100100000011:	sigmoid = 21'b111111111111111111000;
		14'b01100100000100:	sigmoid = 21'b111111111111111111000;
		14'b01100100000101:	sigmoid = 21'b111111111111111111000;
		14'b01100100000110:	sigmoid = 21'b111111111111111111000;
		14'b01100100000111:	sigmoid = 21'b111111111111111111000;
		14'b01100100001000:	sigmoid = 21'b111111111111111111000;
		14'b01100100001001:	sigmoid = 21'b111111111111111111000;
		14'b01100100001010:	sigmoid = 21'b111111111111111111000;
		14'b01100100001011:	sigmoid = 21'b111111111111111111000;
		14'b01100100001100:	sigmoid = 21'b111111111111111111000;
		14'b01100100001101:	sigmoid = 21'b111111111111111111000;
		14'b01100100001110:	sigmoid = 21'b111111111111111111000;
		14'b01100100001111:	sigmoid = 21'b111111111111111111000;
		14'b01100100010000:	sigmoid = 21'b111111111111111111000;
		14'b01100100010001:	sigmoid = 21'b111111111111111111000;
		14'b01100100010010:	sigmoid = 21'b111111111111111111000;
		14'b01100100010011:	sigmoid = 21'b111111111111111111000;
		14'b01100100010100:	sigmoid = 21'b111111111111111111000;
		14'b01100100010101:	sigmoid = 21'b111111111111111111000;
		14'b01100100010110:	sigmoid = 21'b111111111111111111000;
		14'b01100100010111:	sigmoid = 21'b111111111111111111000;
		14'b01100100011000:	sigmoid = 21'b111111111111111111000;
		14'b01100100011001:	sigmoid = 21'b111111111111111111000;
		14'b01100100011010:	sigmoid = 21'b111111111111111111000;
		14'b01100100011011:	sigmoid = 21'b111111111111111111000;
		14'b01100100011100:	sigmoid = 21'b111111111111111111000;
		14'b01100100011101:	sigmoid = 21'b111111111111111111000;
		14'b01100100011110:	sigmoid = 21'b111111111111111111000;
		14'b01100100011111:	sigmoid = 21'b111111111111111111000;
		14'b01100100100000:	sigmoid = 21'b111111111111111111000;
		14'b01100100100001:	sigmoid = 21'b111111111111111111000;
		14'b01100100100010:	sigmoid = 21'b111111111111111111000;
		14'b01100100100011:	sigmoid = 21'b111111111111111111000;
		14'b01100100100100:	sigmoid = 21'b111111111111111111000;
		14'b01100100100101:	sigmoid = 21'b111111111111111111000;
		14'b01100100100110:	sigmoid = 21'b111111111111111111000;
		14'b01100100100111:	sigmoid = 21'b111111111111111111000;
		14'b01100100101000:	sigmoid = 21'b111111111111111111000;
		14'b01100100101001:	sigmoid = 21'b111111111111111111000;
		14'b01100100101010:	sigmoid = 21'b111111111111111111000;
		14'b01100100101011:	sigmoid = 21'b111111111111111111000;
		14'b01100100101100:	sigmoid = 21'b111111111111111111000;
		14'b01100100101101:	sigmoid = 21'b111111111111111111000;
		14'b01100100101110:	sigmoid = 21'b111111111111111111000;
		14'b01100100101111:	sigmoid = 21'b111111111111111111000;
		14'b01100100110000:	sigmoid = 21'b111111111111111111000;
		14'b01100100110001:	sigmoid = 21'b111111111111111111000;
		14'b01100100110010:	sigmoid = 21'b111111111111111111000;
		14'b01100100110011:	sigmoid = 21'b111111111111111111000;
		14'b01100100110100:	sigmoid = 21'b111111111111111111000;
		14'b01100100110101:	sigmoid = 21'b111111111111111111000;
		14'b01100100110110:	sigmoid = 21'b111111111111111111000;
		14'b01100100110111:	sigmoid = 21'b111111111111111111000;
		14'b01100100111000:	sigmoid = 21'b111111111111111111000;
		14'b01100100111001:	sigmoid = 21'b111111111111111111001;
		14'b01100100111010:	sigmoid = 21'b111111111111111111001;
		14'b01100100111011:	sigmoid = 21'b111111111111111111001;
		14'b01100100111100:	sigmoid = 21'b111111111111111111001;
		14'b01100100111101:	sigmoid = 21'b111111111111111111001;
		14'b01100100111110:	sigmoid = 21'b111111111111111111001;
		14'b01100100111111:	sigmoid = 21'b111111111111111111001;
		14'b01100101000000:	sigmoid = 21'b111111111111111111001;
		14'b01100101000001:	sigmoid = 21'b111111111111111111001;
		14'b01100101000010:	sigmoid = 21'b111111111111111111001;
		14'b01100101000011:	sigmoid = 21'b111111111111111111001;
		14'b01100101000100:	sigmoid = 21'b111111111111111111001;
		14'b01100101000101:	sigmoid = 21'b111111111111111111001;
		14'b01100101000110:	sigmoid = 21'b111111111111111111001;
		14'b01100101000111:	sigmoid = 21'b111111111111111111001;
		14'b01100101001000:	sigmoid = 21'b111111111111111111001;
		14'b01100101001001:	sigmoid = 21'b111111111111111111001;
		14'b01100101001010:	sigmoid = 21'b111111111111111111001;
		14'b01100101001011:	sigmoid = 21'b111111111111111111001;
		14'b01100101001100:	sigmoid = 21'b111111111111111111001;
		14'b01100101001101:	sigmoid = 21'b111111111111111111001;
		14'b01100101001110:	sigmoid = 21'b111111111111111111001;
		14'b01100101001111:	sigmoid = 21'b111111111111111111001;
		14'b01100101010000:	sigmoid = 21'b111111111111111111001;
		14'b01100101010001:	sigmoid = 21'b111111111111111111001;
		14'b01100101010010:	sigmoid = 21'b111111111111111111001;
		14'b01100101010011:	sigmoid = 21'b111111111111111111001;
		14'b01100101010100:	sigmoid = 21'b111111111111111111001;
		14'b01100101010101:	sigmoid = 21'b111111111111111111001;
		14'b01100101010110:	sigmoid = 21'b111111111111111111001;
		14'b01100101010111:	sigmoid = 21'b111111111111111111001;
		14'b01100101011000:	sigmoid = 21'b111111111111111111001;
		14'b01100101011001:	sigmoid = 21'b111111111111111111001;
		14'b01100101011010:	sigmoid = 21'b111111111111111111001;
		14'b01100101011011:	sigmoid = 21'b111111111111111111001;
		14'b01100101011100:	sigmoid = 21'b111111111111111111001;
		14'b01100101011101:	sigmoid = 21'b111111111111111111001;
		14'b01100101011110:	sigmoid = 21'b111111111111111111001;
		14'b01100101011111:	sigmoid = 21'b111111111111111111001;
		14'b01100101100000:	sigmoid = 21'b111111111111111111001;
		14'b01100101100001:	sigmoid = 21'b111111111111111111001;
		14'b01100101100010:	sigmoid = 21'b111111111111111111001;
		14'b01100101100011:	sigmoid = 21'b111111111111111111001;
		14'b01100101100100:	sigmoid = 21'b111111111111111111001;
		14'b01100101100101:	sigmoid = 21'b111111111111111111001;
		14'b01100101100110:	sigmoid = 21'b111111111111111111001;
		14'b01100101100111:	sigmoid = 21'b111111111111111111001;
		14'b01100101101000:	sigmoid = 21'b111111111111111111001;
		14'b01100101101001:	sigmoid = 21'b111111111111111111001;
		14'b01100101101010:	sigmoid = 21'b111111111111111111001;
		14'b01100101101011:	sigmoid = 21'b111111111111111111001;
		14'b01100101101100:	sigmoid = 21'b111111111111111111001;
		14'b01100101101101:	sigmoid = 21'b111111111111111111001;
		14'b01100101101110:	sigmoid = 21'b111111111111111111001;
		14'b01100101101111:	sigmoid = 21'b111111111111111111001;
		14'b01100101110000:	sigmoid = 21'b111111111111111111001;
		14'b01100101110001:	sigmoid = 21'b111111111111111111001;
		14'b01100101110010:	sigmoid = 21'b111111111111111111001;
		14'b01100101110011:	sigmoid = 21'b111111111111111111001;
		14'b01100101110100:	sigmoid = 21'b111111111111111111001;
		14'b01100101110101:	sigmoid = 21'b111111111111111111001;
		14'b01100101110110:	sigmoid = 21'b111111111111111111001;
		14'b01100101110111:	sigmoid = 21'b111111111111111111001;
		14'b01100101111000:	sigmoid = 21'b111111111111111111001;
		14'b01100101111001:	sigmoid = 21'b111111111111111111001;
		14'b01100101111010:	sigmoid = 21'b111111111111111111001;
		14'b01100101111011:	sigmoid = 21'b111111111111111111001;
		14'b01100101111100:	sigmoid = 21'b111111111111111111001;
		14'b01100101111101:	sigmoid = 21'b111111111111111111001;
		14'b01100101111110:	sigmoid = 21'b111111111111111111001;
		14'b01100101111111:	sigmoid = 21'b111111111111111111001;
		14'b01100110000000:	sigmoid = 21'b111111111111111111001;
		14'b01100110000001:	sigmoid = 21'b111111111111111111001;
		14'b01100110000010:	sigmoid = 21'b111111111111111111001;
		14'b01100110000011:	sigmoid = 21'b111111111111111111001;
		14'b01100110000100:	sigmoid = 21'b111111111111111111001;
		14'b01100110000101:	sigmoid = 21'b111111111111111111001;
		14'b01100110000110:	sigmoid = 21'b111111111111111111001;
		14'b01100110000111:	sigmoid = 21'b111111111111111111001;
		14'b01100110001000:	sigmoid = 21'b111111111111111111010;
		14'b01100110001001:	sigmoid = 21'b111111111111111111010;
		14'b01100110001010:	sigmoid = 21'b111111111111111111010;
		14'b01100110001011:	sigmoid = 21'b111111111111111111010;
		14'b01100110001100:	sigmoid = 21'b111111111111111111010;
		14'b01100110001101:	sigmoid = 21'b111111111111111111010;
		14'b01100110001110:	sigmoid = 21'b111111111111111111010;
		14'b01100110001111:	sigmoid = 21'b111111111111111111010;
		14'b01100110010000:	sigmoid = 21'b111111111111111111010;
		14'b01100110010001:	sigmoid = 21'b111111111111111111010;
		14'b01100110010010:	sigmoid = 21'b111111111111111111010;
		14'b01100110010011:	sigmoid = 21'b111111111111111111010;
		14'b01100110010100:	sigmoid = 21'b111111111111111111010;
		14'b01100110010101:	sigmoid = 21'b111111111111111111010;
		14'b01100110010110:	sigmoid = 21'b111111111111111111010;
		14'b01100110010111:	sigmoid = 21'b111111111111111111010;
		14'b01100110011000:	sigmoid = 21'b111111111111111111010;
		14'b01100110011001:	sigmoid = 21'b111111111111111111010;
		14'b01100110011010:	sigmoid = 21'b111111111111111111010;
		14'b01100110011011:	sigmoid = 21'b111111111111111111010;
		14'b01100110011100:	sigmoid = 21'b111111111111111111010;
		14'b01100110011101:	sigmoid = 21'b111111111111111111010;
		14'b01100110011110:	sigmoid = 21'b111111111111111111010;
		14'b01100110011111:	sigmoid = 21'b111111111111111111010;
		14'b01100110100000:	sigmoid = 21'b111111111111111111010;
		14'b01100110100001:	sigmoid = 21'b111111111111111111010;
		14'b01100110100010:	sigmoid = 21'b111111111111111111010;
		14'b01100110100011:	sigmoid = 21'b111111111111111111010;
		14'b01100110100100:	sigmoid = 21'b111111111111111111010;
		14'b01100110100101:	sigmoid = 21'b111111111111111111010;
		14'b01100110100110:	sigmoid = 21'b111111111111111111010;
		14'b01100110100111:	sigmoid = 21'b111111111111111111010;
		14'b01100110101000:	sigmoid = 21'b111111111111111111010;
		14'b01100110101001:	sigmoid = 21'b111111111111111111010;
		14'b01100110101010:	sigmoid = 21'b111111111111111111010;
		14'b01100110101011:	sigmoid = 21'b111111111111111111010;
		14'b01100110101100:	sigmoid = 21'b111111111111111111010;
		14'b01100110101101:	sigmoid = 21'b111111111111111111010;
		14'b01100110101110:	sigmoid = 21'b111111111111111111010;
		14'b01100110101111:	sigmoid = 21'b111111111111111111010;
		14'b01100110110000:	sigmoid = 21'b111111111111111111010;
		14'b01100110110001:	sigmoid = 21'b111111111111111111010;
		14'b01100110110010:	sigmoid = 21'b111111111111111111010;
		14'b01100110110011:	sigmoid = 21'b111111111111111111010;
		14'b01100110110100:	sigmoid = 21'b111111111111111111010;
		14'b01100110110101:	sigmoid = 21'b111111111111111111010;
		14'b01100110110110:	sigmoid = 21'b111111111111111111010;
		14'b01100110110111:	sigmoid = 21'b111111111111111111010;
		14'b01100110111000:	sigmoid = 21'b111111111111111111010;
		14'b01100110111001:	sigmoid = 21'b111111111111111111010;
		14'b01100110111010:	sigmoid = 21'b111111111111111111010;
		14'b01100110111011:	sigmoid = 21'b111111111111111111010;
		14'b01100110111100:	sigmoid = 21'b111111111111111111010;
		14'b01100110111101:	sigmoid = 21'b111111111111111111010;
		14'b01100110111110:	sigmoid = 21'b111111111111111111010;
		14'b01100110111111:	sigmoid = 21'b111111111111111111010;
		14'b01100111000000:	sigmoid = 21'b111111111111111111010;
		14'b01100111000001:	sigmoid = 21'b111111111111111111010;
		14'b01100111000010:	sigmoid = 21'b111111111111111111010;
		14'b01100111000011:	sigmoid = 21'b111111111111111111010;
		14'b01100111000100:	sigmoid = 21'b111111111111111111010;
		14'b01100111000101:	sigmoid = 21'b111111111111111111010;
		14'b01100111000110:	sigmoid = 21'b111111111111111111010;
		14'b01100111000111:	sigmoid = 21'b111111111111111111010;
		14'b01100111001000:	sigmoid = 21'b111111111111111111010;
		14'b01100111001001:	sigmoid = 21'b111111111111111111010;
		14'b01100111001010:	sigmoid = 21'b111111111111111111010;
		14'b01100111001011:	sigmoid = 21'b111111111111111111010;
		14'b01100111001100:	sigmoid = 21'b111111111111111111010;
		14'b01100111001101:	sigmoid = 21'b111111111111111111010;
		14'b01100111001110:	sigmoid = 21'b111111111111111111010;
		14'b01100111001111:	sigmoid = 21'b111111111111111111010;
		14'b01100111010000:	sigmoid = 21'b111111111111111111010;
		14'b01100111010001:	sigmoid = 21'b111111111111111111010;
		14'b01100111010010:	sigmoid = 21'b111111111111111111010;
		14'b01100111010011:	sigmoid = 21'b111111111111111111010;
		14'b01100111010100:	sigmoid = 21'b111111111111111111010;
		14'b01100111010101:	sigmoid = 21'b111111111111111111010;
		14'b01100111010110:	sigmoid = 21'b111111111111111111010;
		14'b01100111010111:	sigmoid = 21'b111111111111111111010;
		14'b01100111011000:	sigmoid = 21'b111111111111111111010;
		14'b01100111011001:	sigmoid = 21'b111111111111111111010;
		14'b01100111011010:	sigmoid = 21'b111111111111111111010;
		14'b01100111011011:	sigmoid = 21'b111111111111111111010;
		14'b01100111011100:	sigmoid = 21'b111111111111111111010;
		14'b01100111011101:	sigmoid = 21'b111111111111111111010;
		14'b01100111011110:	sigmoid = 21'b111111111111111111010;
		14'b01100111011111:	sigmoid = 21'b111111111111111111010;
		14'b01100111100000:	sigmoid = 21'b111111111111111111010;
		14'b01100111100001:	sigmoid = 21'b111111111111111111010;
		14'b01100111100010:	sigmoid = 21'b111111111111111111010;
		14'b01100111100011:	sigmoid = 21'b111111111111111111010;
		14'b01100111100100:	sigmoid = 21'b111111111111111111010;
		14'b01100111100101:	sigmoid = 21'b111111111111111111011;
		14'b01100111100110:	sigmoid = 21'b111111111111111111011;
		14'b01100111100111:	sigmoid = 21'b111111111111111111011;
		14'b01100111101000:	sigmoid = 21'b111111111111111111011;
		14'b01100111101001:	sigmoid = 21'b111111111111111111011;
		14'b01100111101010:	sigmoid = 21'b111111111111111111011;
		14'b01100111101011:	sigmoid = 21'b111111111111111111011;
		14'b01100111101100:	sigmoid = 21'b111111111111111111011;
		14'b01100111101101:	sigmoid = 21'b111111111111111111011;
		14'b01100111101110:	sigmoid = 21'b111111111111111111011;
		14'b01100111101111:	sigmoid = 21'b111111111111111111011;
		14'b01100111110000:	sigmoid = 21'b111111111111111111011;
		14'b01100111110001:	sigmoid = 21'b111111111111111111011;
		14'b01100111110010:	sigmoid = 21'b111111111111111111011;
		14'b01100111110011:	sigmoid = 21'b111111111111111111011;
		14'b01100111110100:	sigmoid = 21'b111111111111111111011;
		14'b01100111110101:	sigmoid = 21'b111111111111111111011;
		14'b01100111110110:	sigmoid = 21'b111111111111111111011;
		14'b01100111110111:	sigmoid = 21'b111111111111111111011;
		14'b01100111111000:	sigmoid = 21'b111111111111111111011;
		14'b01100111111001:	sigmoid = 21'b111111111111111111011;
		14'b01100111111010:	sigmoid = 21'b111111111111111111011;
		14'b01100111111011:	sigmoid = 21'b111111111111111111011;
		14'b01100111111100:	sigmoid = 21'b111111111111111111011;
		14'b01100111111101:	sigmoid = 21'b111111111111111111011;
		14'b01100111111110:	sigmoid = 21'b111111111111111111011;
		14'b01100111111111:	sigmoid = 21'b111111111111111111011;
		14'b01101000000000:	sigmoid = 21'b111111111111111111011;
		14'b01101000000001:	sigmoid = 21'b111111111111111111011;
		14'b01101000000010:	sigmoid = 21'b111111111111111111011;
		14'b01101000000011:	sigmoid = 21'b111111111111111111011;
		14'b01101000000100:	sigmoid = 21'b111111111111111111011;
		14'b01101000000101:	sigmoid = 21'b111111111111111111011;
		14'b01101000000110:	sigmoid = 21'b111111111111111111011;
		14'b01101000000111:	sigmoid = 21'b111111111111111111011;
		14'b01101000001000:	sigmoid = 21'b111111111111111111011;
		14'b01101000001001:	sigmoid = 21'b111111111111111111011;
		14'b01101000001010:	sigmoid = 21'b111111111111111111011;
		14'b01101000001011:	sigmoid = 21'b111111111111111111011;
		14'b01101000001100:	sigmoid = 21'b111111111111111111011;
		14'b01101000001101:	sigmoid = 21'b111111111111111111011;
		14'b01101000001110:	sigmoid = 21'b111111111111111111011;
		14'b01101000001111:	sigmoid = 21'b111111111111111111011;
		14'b01101000010000:	sigmoid = 21'b111111111111111111011;
		14'b01101000010001:	sigmoid = 21'b111111111111111111011;
		14'b01101000010010:	sigmoid = 21'b111111111111111111011;
		14'b01101000010011:	sigmoid = 21'b111111111111111111011;
		14'b01101000010100:	sigmoid = 21'b111111111111111111011;
		14'b01101000010101:	sigmoid = 21'b111111111111111111011;
		14'b01101000010110:	sigmoid = 21'b111111111111111111011;
		14'b01101000010111:	sigmoid = 21'b111111111111111111011;
		14'b01101000011000:	sigmoid = 21'b111111111111111111011;
		14'b01101000011001:	sigmoid = 21'b111111111111111111011;
		14'b01101000011010:	sigmoid = 21'b111111111111111111011;
		14'b01101000011011:	sigmoid = 21'b111111111111111111011;
		14'b01101000011100:	sigmoid = 21'b111111111111111111011;
		14'b01101000011101:	sigmoid = 21'b111111111111111111011;
		14'b01101000011110:	sigmoid = 21'b111111111111111111011;
		14'b01101000011111:	sigmoid = 21'b111111111111111111011;
		14'b01101000100000:	sigmoid = 21'b111111111111111111011;
		14'b01101000100001:	sigmoid = 21'b111111111111111111011;
		14'b01101000100010:	sigmoid = 21'b111111111111111111011;
		14'b01101000100011:	sigmoid = 21'b111111111111111111011;
		14'b01101000100100:	sigmoid = 21'b111111111111111111011;
		14'b01101000100101:	sigmoid = 21'b111111111111111111011;
		14'b01101000100110:	sigmoid = 21'b111111111111111111011;
		14'b01101000100111:	sigmoid = 21'b111111111111111111011;
		14'b01101000101000:	sigmoid = 21'b111111111111111111011;
		14'b01101000101001:	sigmoid = 21'b111111111111111111011;
		14'b01101000101010:	sigmoid = 21'b111111111111111111011;
		14'b01101000101011:	sigmoid = 21'b111111111111111111011;
		14'b01101000101100:	sigmoid = 21'b111111111111111111011;
		14'b01101000101101:	sigmoid = 21'b111111111111111111011;
		14'b01101000101110:	sigmoid = 21'b111111111111111111011;
		14'b01101000101111:	sigmoid = 21'b111111111111111111011;
		14'b01101000110000:	sigmoid = 21'b111111111111111111011;
		14'b01101000110001:	sigmoid = 21'b111111111111111111011;
		14'b01101000110010:	sigmoid = 21'b111111111111111111011;
		14'b01101000110011:	sigmoid = 21'b111111111111111111011;
		14'b01101000110100:	sigmoid = 21'b111111111111111111011;
		14'b01101000110101:	sigmoid = 21'b111111111111111111011;
		14'b01101000110110:	sigmoid = 21'b111111111111111111011;
		14'b01101000110111:	sigmoid = 21'b111111111111111111011;
		14'b01101000111000:	sigmoid = 21'b111111111111111111011;
		14'b01101000111001:	sigmoid = 21'b111111111111111111011;
		14'b01101000111010:	sigmoid = 21'b111111111111111111011;
		14'b01101000111011:	sigmoid = 21'b111111111111111111011;
		14'b01101000111100:	sigmoid = 21'b111111111111111111011;
		14'b01101000111101:	sigmoid = 21'b111111111111111111011;
		14'b01101000111110:	sigmoid = 21'b111111111111111111011;
		14'b01101000111111:	sigmoid = 21'b111111111111111111011;
		14'b01101001000000:	sigmoid = 21'b111111111111111111011;
		14'b01101001000001:	sigmoid = 21'b111111111111111111011;
		14'b01101001000010:	sigmoid = 21'b111111111111111111011;
		14'b01101001000011:	sigmoid = 21'b111111111111111111011;
		14'b01101001000100:	sigmoid = 21'b111111111111111111011;
		14'b01101001000101:	sigmoid = 21'b111111111111111111011;
		14'b01101001000110:	sigmoid = 21'b111111111111111111011;
		14'b01101001000111:	sigmoid = 21'b111111111111111111011;
		14'b01101001001000:	sigmoid = 21'b111111111111111111011;
		14'b01101001001001:	sigmoid = 21'b111111111111111111011;
		14'b01101001001010:	sigmoid = 21'b111111111111111111011;
		14'b01101001001011:	sigmoid = 21'b111111111111111111011;
		14'b01101001001100:	sigmoid = 21'b111111111111111111011;
		14'b01101001001101:	sigmoid = 21'b111111111111111111011;
		14'b01101001001110:	sigmoid = 21'b111111111111111111011;
		14'b01101001001111:	sigmoid = 21'b111111111111111111011;
		14'b01101001010000:	sigmoid = 21'b111111111111111111011;
		14'b01101001010001:	sigmoid = 21'b111111111111111111011;
		14'b01101001010010:	sigmoid = 21'b111111111111111111011;
		14'b01101001010011:	sigmoid = 21'b111111111111111111011;
		14'b01101001010100:	sigmoid = 21'b111111111111111111011;
		14'b01101001010101:	sigmoid = 21'b111111111111111111011;
		14'b01101001010110:	sigmoid = 21'b111111111111111111011;
		14'b01101001010111:	sigmoid = 21'b111111111111111111100;
		14'b01101001011000:	sigmoid = 21'b111111111111111111100;
		14'b01101001011001:	sigmoid = 21'b111111111111111111100;
		14'b01101001011010:	sigmoid = 21'b111111111111111111100;
		14'b01101001011011:	sigmoid = 21'b111111111111111111100;
		14'b01101001011100:	sigmoid = 21'b111111111111111111100;
		14'b01101001011101:	sigmoid = 21'b111111111111111111100;
		14'b01101001011110:	sigmoid = 21'b111111111111111111100;
		14'b01101001011111:	sigmoid = 21'b111111111111111111100;
		14'b01101001100000:	sigmoid = 21'b111111111111111111100;
		14'b01101001100001:	sigmoid = 21'b111111111111111111100;
		14'b01101001100010:	sigmoid = 21'b111111111111111111100;
		14'b01101001100011:	sigmoid = 21'b111111111111111111100;
		14'b01101001100100:	sigmoid = 21'b111111111111111111100;
		14'b01101001100101:	sigmoid = 21'b111111111111111111100;
		14'b01101001100110:	sigmoid = 21'b111111111111111111100;
		14'b01101001100111:	sigmoid = 21'b111111111111111111100;
		14'b01101001101000:	sigmoid = 21'b111111111111111111100;
		14'b01101001101001:	sigmoid = 21'b111111111111111111100;
		14'b01101001101010:	sigmoid = 21'b111111111111111111100;
		14'b01101001101011:	sigmoid = 21'b111111111111111111100;
		14'b01101001101100:	sigmoid = 21'b111111111111111111100;
		14'b01101001101101:	sigmoid = 21'b111111111111111111100;
		14'b01101001101110:	sigmoid = 21'b111111111111111111100;
		14'b01101001101111:	sigmoid = 21'b111111111111111111100;
		14'b01101001110000:	sigmoid = 21'b111111111111111111100;
		14'b01101001110001:	sigmoid = 21'b111111111111111111100;
		14'b01101001110010:	sigmoid = 21'b111111111111111111100;
		14'b01101001110011:	sigmoid = 21'b111111111111111111100;
		14'b01101001110100:	sigmoid = 21'b111111111111111111100;
		14'b01101001110101:	sigmoid = 21'b111111111111111111100;
		14'b01101001110110:	sigmoid = 21'b111111111111111111100;
		14'b01101001110111:	sigmoid = 21'b111111111111111111100;
		14'b01101001111000:	sigmoid = 21'b111111111111111111100;
		14'b01101001111001:	sigmoid = 21'b111111111111111111100;
		14'b01101001111010:	sigmoid = 21'b111111111111111111100;
		14'b01101001111011:	sigmoid = 21'b111111111111111111100;
		14'b01101001111100:	sigmoid = 21'b111111111111111111100;
		14'b01101001111101:	sigmoid = 21'b111111111111111111100;
		14'b01101001111110:	sigmoid = 21'b111111111111111111100;
		14'b01101001111111:	sigmoid = 21'b111111111111111111100;
		14'b01101010000000:	sigmoid = 21'b111111111111111111100;
		14'b01101010000001:	sigmoid = 21'b111111111111111111100;
		14'b01101010000010:	sigmoid = 21'b111111111111111111100;
		14'b01101010000011:	sigmoid = 21'b111111111111111111100;
		14'b01101010000100:	sigmoid = 21'b111111111111111111100;
		14'b01101010000101:	sigmoid = 21'b111111111111111111100;
		14'b01101010000110:	sigmoid = 21'b111111111111111111100;
		14'b01101010000111:	sigmoid = 21'b111111111111111111100;
		14'b01101010001000:	sigmoid = 21'b111111111111111111100;
		14'b01101010001001:	sigmoid = 21'b111111111111111111100;
		14'b01101010001010:	sigmoid = 21'b111111111111111111100;
		14'b01101010001011:	sigmoid = 21'b111111111111111111100;
		14'b01101010001100:	sigmoid = 21'b111111111111111111100;
		14'b01101010001101:	sigmoid = 21'b111111111111111111100;
		14'b01101010001110:	sigmoid = 21'b111111111111111111100;
		14'b01101010001111:	sigmoid = 21'b111111111111111111100;
		14'b01101010010000:	sigmoid = 21'b111111111111111111100;
		14'b01101010010001:	sigmoid = 21'b111111111111111111100;
		14'b01101010010010:	sigmoid = 21'b111111111111111111100;
		14'b01101010010011:	sigmoid = 21'b111111111111111111100;
		14'b01101010010100:	sigmoid = 21'b111111111111111111100;
		14'b01101010010101:	sigmoid = 21'b111111111111111111100;
		14'b01101010010110:	sigmoid = 21'b111111111111111111100;
		14'b01101010010111:	sigmoid = 21'b111111111111111111100;
		14'b01101010011000:	sigmoid = 21'b111111111111111111100;
		14'b01101010011001:	sigmoid = 21'b111111111111111111100;
		14'b01101010011010:	sigmoid = 21'b111111111111111111100;
		14'b01101010011011:	sigmoid = 21'b111111111111111111100;
		14'b01101010011100:	sigmoid = 21'b111111111111111111100;
		14'b01101010011101:	sigmoid = 21'b111111111111111111100;
		14'b01101010011110:	sigmoid = 21'b111111111111111111100;
		14'b01101010011111:	sigmoid = 21'b111111111111111111100;
		14'b01101010100000:	sigmoid = 21'b111111111111111111100;
		14'b01101010100001:	sigmoid = 21'b111111111111111111100;
		14'b01101010100010:	sigmoid = 21'b111111111111111111100;
		14'b01101010100011:	sigmoid = 21'b111111111111111111100;
		14'b01101010100100:	sigmoid = 21'b111111111111111111100;
		14'b01101010100101:	sigmoid = 21'b111111111111111111100;
		14'b01101010100110:	sigmoid = 21'b111111111111111111100;
		14'b01101010100111:	sigmoid = 21'b111111111111111111100;
		14'b01101010101000:	sigmoid = 21'b111111111111111111100;
		14'b01101010101001:	sigmoid = 21'b111111111111111111100;
		14'b01101010101010:	sigmoid = 21'b111111111111111111100;
		14'b01101010101011:	sigmoid = 21'b111111111111111111100;
		14'b01101010101100:	sigmoid = 21'b111111111111111111100;
		14'b01101010101101:	sigmoid = 21'b111111111111111111100;
		14'b01101010101110:	sigmoid = 21'b111111111111111111100;
		14'b01101010101111:	sigmoid = 21'b111111111111111111100;
		14'b01101010110000:	sigmoid = 21'b111111111111111111100;
		14'b01101010110001:	sigmoid = 21'b111111111111111111100;
		14'b01101010110010:	sigmoid = 21'b111111111111111111100;
		14'b01101010110011:	sigmoid = 21'b111111111111111111100;
		14'b01101010110100:	sigmoid = 21'b111111111111111111100;
		14'b01101010110101:	sigmoid = 21'b111111111111111111100;
		14'b01101010110110:	sigmoid = 21'b111111111111111111100;
		14'b01101010110111:	sigmoid = 21'b111111111111111111100;
		14'b01101010111000:	sigmoid = 21'b111111111111111111100;
		14'b01101010111001:	sigmoid = 21'b111111111111111111100;
		14'b01101010111010:	sigmoid = 21'b111111111111111111100;
		14'b01101010111011:	sigmoid = 21'b111111111111111111100;
		14'b01101010111100:	sigmoid = 21'b111111111111111111100;
		14'b01101010111101:	sigmoid = 21'b111111111111111111100;
		14'b01101010111110:	sigmoid = 21'b111111111111111111100;
		14'b01101010111111:	sigmoid = 21'b111111111111111111100;
		14'b01101011000000:	sigmoid = 21'b111111111111111111100;
		14'b01101011000001:	sigmoid = 21'b111111111111111111100;
		14'b01101011000010:	sigmoid = 21'b111111111111111111100;
		14'b01101011000011:	sigmoid = 21'b111111111111111111100;
		14'b01101011000100:	sigmoid = 21'b111111111111111111100;
		14'b01101011000101:	sigmoid = 21'b111111111111111111100;
		14'b01101011000110:	sigmoid = 21'b111111111111111111100;
		14'b01101011000111:	sigmoid = 21'b111111111111111111100;
		14'b01101011001000:	sigmoid = 21'b111111111111111111100;
		14'b01101011001001:	sigmoid = 21'b111111111111111111100;
		14'b01101011001010:	sigmoid = 21'b111111111111111111100;
		14'b01101011001011:	sigmoid = 21'b111111111111111111100;
		14'b01101011001100:	sigmoid = 21'b111111111111111111100;
		14'b01101011001101:	sigmoid = 21'b111111111111111111100;
		14'b01101011001110:	sigmoid = 21'b111111111111111111100;
		14'b01101011001111:	sigmoid = 21'b111111111111111111100;
		14'b01101011010000:	sigmoid = 21'b111111111111111111100;
		14'b01101011010001:	sigmoid = 21'b111111111111111111100;
		14'b01101011010010:	sigmoid = 21'b111111111111111111100;
		14'b01101011010011:	sigmoid = 21'b111111111111111111100;
		14'b01101011010100:	sigmoid = 21'b111111111111111111100;
		14'b01101011010101:	sigmoid = 21'b111111111111111111100;
		14'b01101011010110:	sigmoid = 21'b111111111111111111100;
		14'b01101011010111:	sigmoid = 21'b111111111111111111100;
		14'b01101011011000:	sigmoid = 21'b111111111111111111100;
		14'b01101011011001:	sigmoid = 21'b111111111111111111100;
		14'b01101011011010:	sigmoid = 21'b111111111111111111100;
		14'b01101011011011:	sigmoid = 21'b111111111111111111100;
		14'b01101011011100:	sigmoid = 21'b111111111111111111100;
		14'b01101011011101:	sigmoid = 21'b111111111111111111100;
		14'b01101011011110:	sigmoid = 21'b111111111111111111100;
		14'b01101011011111:	sigmoid = 21'b111111111111111111100;
		14'b01101011100000:	sigmoid = 21'b111111111111111111100;
		14'b01101011100001:	sigmoid = 21'b111111111111111111100;
		14'b01101011100010:	sigmoid = 21'b111111111111111111100;
		14'b01101011100011:	sigmoid = 21'b111111111111111111100;
		14'b01101011100100:	sigmoid = 21'b111111111111111111100;
		14'b01101011100101:	sigmoid = 21'b111111111111111111100;
		14'b01101011100110:	sigmoid = 21'b111111111111111111100;
		14'b01101011100111:	sigmoid = 21'b111111111111111111100;
		14'b01101011101000:	sigmoid = 21'b111111111111111111100;
		14'b01101011101001:	sigmoid = 21'b111111111111111111100;
		14'b01101011101010:	sigmoid = 21'b111111111111111111100;
		14'b01101011101011:	sigmoid = 21'b111111111111111111101;
		14'b01101011101100:	sigmoid = 21'b111111111111111111101;
		14'b01101011101101:	sigmoid = 21'b111111111111111111101;
		14'b01101011101110:	sigmoid = 21'b111111111111111111101;
		14'b01101011101111:	sigmoid = 21'b111111111111111111101;
		14'b01101011110000:	sigmoid = 21'b111111111111111111101;
		14'b01101011110001:	sigmoid = 21'b111111111111111111101;
		14'b01101011110010:	sigmoid = 21'b111111111111111111101;
		14'b01101011110011:	sigmoid = 21'b111111111111111111101;
		14'b01101011110100:	sigmoid = 21'b111111111111111111101;
		14'b01101011110101:	sigmoid = 21'b111111111111111111101;
		14'b01101011110110:	sigmoid = 21'b111111111111111111101;
		14'b01101011110111:	sigmoid = 21'b111111111111111111101;
		14'b01101011111000:	sigmoid = 21'b111111111111111111101;
		14'b01101011111001:	sigmoid = 21'b111111111111111111101;
		14'b01101011111010:	sigmoid = 21'b111111111111111111101;
		14'b01101011111011:	sigmoid = 21'b111111111111111111101;
		14'b01101011111100:	sigmoid = 21'b111111111111111111101;
		14'b01101011111101:	sigmoid = 21'b111111111111111111101;
		14'b01101011111110:	sigmoid = 21'b111111111111111111101;
		14'b01101011111111:	sigmoid = 21'b111111111111111111101;
		14'b01101100000000:	sigmoid = 21'b111111111111111111101;
		14'b01101100000001:	sigmoid = 21'b111111111111111111101;
		14'b01101100000010:	sigmoid = 21'b111111111111111111101;
		14'b01101100000011:	sigmoid = 21'b111111111111111111101;
		14'b01101100000100:	sigmoid = 21'b111111111111111111101;
		14'b01101100000101:	sigmoid = 21'b111111111111111111101;
		14'b01101100000110:	sigmoid = 21'b111111111111111111101;
		14'b01101100000111:	sigmoid = 21'b111111111111111111101;
		14'b01101100001000:	sigmoid = 21'b111111111111111111101;
		14'b01101100001001:	sigmoid = 21'b111111111111111111101;
		14'b01101100001010:	sigmoid = 21'b111111111111111111101;
		14'b01101100001011:	sigmoid = 21'b111111111111111111101;
		14'b01101100001100:	sigmoid = 21'b111111111111111111101;
		14'b01101100001101:	sigmoid = 21'b111111111111111111101;
		14'b01101100001110:	sigmoid = 21'b111111111111111111101;
		14'b01101100001111:	sigmoid = 21'b111111111111111111101;
		14'b01101100010000:	sigmoid = 21'b111111111111111111101;
		14'b01101100010001:	sigmoid = 21'b111111111111111111101;
		14'b01101100010010:	sigmoid = 21'b111111111111111111101;
		14'b01101100010011:	sigmoid = 21'b111111111111111111101;
		14'b01101100010100:	sigmoid = 21'b111111111111111111101;
		14'b01101100010101:	sigmoid = 21'b111111111111111111101;
		14'b01101100010110:	sigmoid = 21'b111111111111111111101;
		14'b01101100010111:	sigmoid = 21'b111111111111111111101;
		14'b01101100011000:	sigmoid = 21'b111111111111111111101;
		14'b01101100011001:	sigmoid = 21'b111111111111111111101;
		14'b01101100011010:	sigmoid = 21'b111111111111111111101;
		14'b01101100011011:	sigmoid = 21'b111111111111111111101;
		14'b01101100011100:	sigmoid = 21'b111111111111111111101;
		14'b01101100011101:	sigmoid = 21'b111111111111111111101;
		14'b01101100011110:	sigmoid = 21'b111111111111111111101;
		14'b01101100011111:	sigmoid = 21'b111111111111111111101;
		14'b01101100100000:	sigmoid = 21'b111111111111111111101;
		14'b01101100100001:	sigmoid = 21'b111111111111111111101;
		14'b01101100100010:	sigmoid = 21'b111111111111111111101;
		14'b01101100100011:	sigmoid = 21'b111111111111111111101;
		14'b01101100100100:	sigmoid = 21'b111111111111111111101;
		14'b01101100100101:	sigmoid = 21'b111111111111111111101;
		14'b01101100100110:	sigmoid = 21'b111111111111111111101;
		14'b01101100100111:	sigmoid = 21'b111111111111111111101;
		14'b01101100101000:	sigmoid = 21'b111111111111111111101;
		14'b01101100101001:	sigmoid = 21'b111111111111111111101;
		14'b01101100101010:	sigmoid = 21'b111111111111111111101;
		14'b01101100101011:	sigmoid = 21'b111111111111111111101;
		14'b01101100101100:	sigmoid = 21'b111111111111111111101;
		14'b01101100101101:	sigmoid = 21'b111111111111111111101;
		14'b01101100101110:	sigmoid = 21'b111111111111111111101;
		14'b01101100101111:	sigmoid = 21'b111111111111111111101;
		14'b01101100110000:	sigmoid = 21'b111111111111111111101;
		14'b01101100110001:	sigmoid = 21'b111111111111111111101;
		14'b01101100110010:	sigmoid = 21'b111111111111111111101;
		14'b01101100110011:	sigmoid = 21'b111111111111111111101;
		14'b01101100110100:	sigmoid = 21'b111111111111111111101;
		14'b01101100110101:	sigmoid = 21'b111111111111111111101;
		14'b01101100110110:	sigmoid = 21'b111111111111111111101;
		14'b01101100110111:	sigmoid = 21'b111111111111111111101;
		14'b01101100111000:	sigmoid = 21'b111111111111111111101;
		14'b01101100111001:	sigmoid = 21'b111111111111111111101;
		14'b01101100111010:	sigmoid = 21'b111111111111111111101;
		14'b01101100111011:	sigmoid = 21'b111111111111111111101;
		14'b01101100111100:	sigmoid = 21'b111111111111111111101;
		14'b01101100111101:	sigmoid = 21'b111111111111111111101;
		14'b01101100111110:	sigmoid = 21'b111111111111111111101;
		14'b01101100111111:	sigmoid = 21'b111111111111111111101;
		14'b01101101000000:	sigmoid = 21'b111111111111111111101;
		14'b01101101000001:	sigmoid = 21'b111111111111111111101;
		14'b01101101000010:	sigmoid = 21'b111111111111111111101;
		14'b01101101000011:	sigmoid = 21'b111111111111111111101;
		14'b01101101000100:	sigmoid = 21'b111111111111111111101;
		14'b01101101000101:	sigmoid = 21'b111111111111111111101;
		14'b01101101000110:	sigmoid = 21'b111111111111111111101;
		14'b01101101000111:	sigmoid = 21'b111111111111111111101;
		14'b01101101001000:	sigmoid = 21'b111111111111111111101;
		14'b01101101001001:	sigmoid = 21'b111111111111111111101;
		14'b01101101001010:	sigmoid = 21'b111111111111111111101;
		14'b01101101001011:	sigmoid = 21'b111111111111111111101;
		14'b01101101001100:	sigmoid = 21'b111111111111111111101;
		14'b01101101001101:	sigmoid = 21'b111111111111111111101;
		14'b01101101001110:	sigmoid = 21'b111111111111111111101;
		14'b01101101001111:	sigmoid = 21'b111111111111111111101;
		14'b01101101010000:	sigmoid = 21'b111111111111111111101;
		14'b01101101010001:	sigmoid = 21'b111111111111111111101;
		14'b01101101010010:	sigmoid = 21'b111111111111111111101;
		14'b01101101010011:	sigmoid = 21'b111111111111111111101;
		14'b01101101010100:	sigmoid = 21'b111111111111111111101;
		14'b01101101010101:	sigmoid = 21'b111111111111111111101;
		14'b01101101010110:	sigmoid = 21'b111111111111111111101;
		14'b01101101010111:	sigmoid = 21'b111111111111111111101;
		14'b01101101011000:	sigmoid = 21'b111111111111111111101;
		14'b01101101011001:	sigmoid = 21'b111111111111111111101;
		14'b01101101011010:	sigmoid = 21'b111111111111111111101;
		14'b01101101011011:	sigmoid = 21'b111111111111111111101;
		14'b01101101011100:	sigmoid = 21'b111111111111111111101;
		14'b01101101011101:	sigmoid = 21'b111111111111111111101;
		14'b01101101011110:	sigmoid = 21'b111111111111111111101;
		14'b01101101011111:	sigmoid = 21'b111111111111111111101;
		14'b01101101100000:	sigmoid = 21'b111111111111111111101;
		14'b01101101100001:	sigmoid = 21'b111111111111111111101;
		14'b01101101100010:	sigmoid = 21'b111111111111111111101;
		14'b01101101100011:	sigmoid = 21'b111111111111111111101;
		14'b01101101100100:	sigmoid = 21'b111111111111111111101;
		14'b01101101100101:	sigmoid = 21'b111111111111111111101;
		14'b01101101100110:	sigmoid = 21'b111111111111111111101;
		14'b01101101100111:	sigmoid = 21'b111111111111111111101;
		14'b01101101101000:	sigmoid = 21'b111111111111111111101;
		14'b01101101101001:	sigmoid = 21'b111111111111111111101;
		14'b01101101101010:	sigmoid = 21'b111111111111111111101;
		14'b01101101101011:	sigmoid = 21'b111111111111111111101;
		14'b01101101101100:	sigmoid = 21'b111111111111111111101;
		14'b01101101101101:	sigmoid = 21'b111111111111111111101;
		14'b01101101101110:	sigmoid = 21'b111111111111111111101;
		14'b01101101101111:	sigmoid = 21'b111111111111111111101;
		14'b01101101110000:	sigmoid = 21'b111111111111111111101;
		14'b01101101110001:	sigmoid = 21'b111111111111111111101;
		14'b01101101110010:	sigmoid = 21'b111111111111111111101;
		14'b01101101110011:	sigmoid = 21'b111111111111111111101;
		14'b01101101110100:	sigmoid = 21'b111111111111111111101;
		14'b01101101110101:	sigmoid = 21'b111111111111111111101;
		14'b01101101110110:	sigmoid = 21'b111111111111111111101;
		14'b01101101110111:	sigmoid = 21'b111111111111111111101;
		14'b01101101111000:	sigmoid = 21'b111111111111111111101;
		14'b01101101111001:	sigmoid = 21'b111111111111111111101;
		14'b01101101111010:	sigmoid = 21'b111111111111111111101;
		14'b01101101111011:	sigmoid = 21'b111111111111111111101;
		14'b01101101111100:	sigmoid = 21'b111111111111111111101;
		14'b01101101111101:	sigmoid = 21'b111111111111111111101;
		14'b01101101111110:	sigmoid = 21'b111111111111111111101;
		14'b01101101111111:	sigmoid = 21'b111111111111111111101;
		14'b01101110000000:	sigmoid = 21'b111111111111111111101;
		14'b01101110000001:	sigmoid = 21'b111111111111111111101;
		14'b01101110000010:	sigmoid = 21'b111111111111111111101;
		14'b01101110000011:	sigmoid = 21'b111111111111111111101;
		14'b01101110000100:	sigmoid = 21'b111111111111111111101;
		14'b01101110000101:	sigmoid = 21'b111111111111111111101;
		14'b01101110000110:	sigmoid = 21'b111111111111111111101;
		14'b01101110000111:	sigmoid = 21'b111111111111111111101;
		14'b01101110001000:	sigmoid = 21'b111111111111111111101;
		14'b01101110001001:	sigmoid = 21'b111111111111111111101;
		14'b01101110001010:	sigmoid = 21'b111111111111111111101;
		14'b01101110001011:	sigmoid = 21'b111111111111111111101;
		14'b01101110001100:	sigmoid = 21'b111111111111111111101;
		14'b01101110001101:	sigmoid = 21'b111111111111111111101;
		14'b01101110001110:	sigmoid = 21'b111111111111111111101;
		14'b01101110001111:	sigmoid = 21'b111111111111111111101;
		14'b01101110010000:	sigmoid = 21'b111111111111111111101;
		14'b01101110010001:	sigmoid = 21'b111111111111111111101;
		14'b01101110010010:	sigmoid = 21'b111111111111111111101;
		14'b01101110010011:	sigmoid = 21'b111111111111111111101;
		14'b01101110010100:	sigmoid = 21'b111111111111111111101;
		14'b01101110010101:	sigmoid = 21'b111111111111111111101;
		14'b01101110010110:	sigmoid = 21'b111111111111111111101;
		14'b01101110010111:	sigmoid = 21'b111111111111111111101;
		14'b01101110011000:	sigmoid = 21'b111111111111111111101;
		14'b01101110011001:	sigmoid = 21'b111111111111111111101;
		14'b01101110011010:	sigmoid = 21'b111111111111111111101;
		14'b01101110011011:	sigmoid = 21'b111111111111111111101;
		14'b01101110011100:	sigmoid = 21'b111111111111111111101;
		14'b01101110011101:	sigmoid = 21'b111111111111111111101;
		14'b01101110011110:	sigmoid = 21'b111111111111111111101;
		14'b01101110011111:	sigmoid = 21'b111111111111111111101;
		14'b01101110100000:	sigmoid = 21'b111111111111111111101;
		14'b01101110100001:	sigmoid = 21'b111111111111111111101;
		14'b01101110100010:	sigmoid = 21'b111111111111111111101;
		14'b01101110100011:	sigmoid = 21'b111111111111111111101;
		14'b01101110100100:	sigmoid = 21'b111111111111111111101;
		14'b01101110100101:	sigmoid = 21'b111111111111111111101;
		14'b01101110100110:	sigmoid = 21'b111111111111111111101;
		14'b01101110100111:	sigmoid = 21'b111111111111111111101;
		14'b01101110101000:	sigmoid = 21'b111111111111111111101;
		14'b01101110101001:	sigmoid = 21'b111111111111111111101;
		14'b01101110101010:	sigmoid = 21'b111111111111111111101;
		14'b01101110101011:	sigmoid = 21'b111111111111111111101;
		14'b01101110101100:	sigmoid = 21'b111111111111111111101;
		14'b01101110101101:	sigmoid = 21'b111111111111111111101;
		14'b01101110101110:	sigmoid = 21'b111111111111111111101;
		14'b01101110101111:	sigmoid = 21'b111111111111111111101;
		14'b01101110110000:	sigmoid = 21'b111111111111111111101;
		14'b01101110110001:	sigmoid = 21'b111111111111111111101;
		14'b01101110110010:	sigmoid = 21'b111111111111111111101;
		14'b01101110110011:	sigmoid = 21'b111111111111111111101;
		14'b01101110110100:	sigmoid = 21'b111111111111111111101;
		14'b01101110110101:	sigmoid = 21'b111111111111111111101;
		14'b01101110110110:	sigmoid = 21'b111111111111111111101;
		14'b01101110110111:	sigmoid = 21'b111111111111111111101;
		14'b01101110111000:	sigmoid = 21'b111111111111111111101;
		14'b01101110111001:	sigmoid = 21'b111111111111111111101;
		14'b01101110111010:	sigmoid = 21'b111111111111111111110;
		14'b01101110111011:	sigmoid = 21'b111111111111111111110;
		14'b01101110111100:	sigmoid = 21'b111111111111111111110;
		14'b01101110111101:	sigmoid = 21'b111111111111111111110;
		14'b01101110111110:	sigmoid = 21'b111111111111111111110;
		14'b01101110111111:	sigmoid = 21'b111111111111111111110;
		14'b01101111000000:	sigmoid = 21'b111111111111111111110;
		14'b01101111000001:	sigmoid = 21'b111111111111111111110;
		14'b01101111000010:	sigmoid = 21'b111111111111111111110;
		14'b01101111000011:	sigmoid = 21'b111111111111111111110;
		14'b01101111000100:	sigmoid = 21'b111111111111111111110;
		14'b01101111000101:	sigmoid = 21'b111111111111111111110;
		14'b01101111000110:	sigmoid = 21'b111111111111111111110;
		14'b01101111000111:	sigmoid = 21'b111111111111111111110;
		14'b01101111001000:	sigmoid = 21'b111111111111111111110;
		14'b01101111001001:	sigmoid = 21'b111111111111111111110;
		14'b01101111001010:	sigmoid = 21'b111111111111111111110;
		14'b01101111001011:	sigmoid = 21'b111111111111111111110;
		14'b01101111001100:	sigmoid = 21'b111111111111111111110;
		14'b01101111001101:	sigmoid = 21'b111111111111111111110;
		14'b01101111001110:	sigmoid = 21'b111111111111111111110;
		14'b01101111001111:	sigmoid = 21'b111111111111111111110;
		14'b01101111010000:	sigmoid = 21'b111111111111111111110;
		14'b01101111010001:	sigmoid = 21'b111111111111111111110;
		14'b01101111010010:	sigmoid = 21'b111111111111111111110;
		14'b01101111010011:	sigmoid = 21'b111111111111111111110;
		14'b01101111010100:	sigmoid = 21'b111111111111111111110;
		14'b01101111010101:	sigmoid = 21'b111111111111111111110;
		14'b01101111010110:	sigmoid = 21'b111111111111111111110;
		14'b01101111010111:	sigmoid = 21'b111111111111111111110;
		14'b01101111011000:	sigmoid = 21'b111111111111111111110;
		14'b01101111011001:	sigmoid = 21'b111111111111111111110;
		14'b01101111011010:	sigmoid = 21'b111111111111111111110;
		14'b01101111011011:	sigmoid = 21'b111111111111111111110;
		14'b01101111011100:	sigmoid = 21'b111111111111111111110;
		14'b01101111011101:	sigmoid = 21'b111111111111111111110;
		14'b01101111011110:	sigmoid = 21'b111111111111111111110;
		14'b01101111011111:	sigmoid = 21'b111111111111111111110;
		14'b01101111100000:	sigmoid = 21'b111111111111111111110;
		14'b01101111100001:	sigmoid = 21'b111111111111111111110;
		14'b01101111100010:	sigmoid = 21'b111111111111111111110;
		14'b01101111100011:	sigmoid = 21'b111111111111111111110;
		14'b01101111100100:	sigmoid = 21'b111111111111111111110;
		14'b01101111100101:	sigmoid = 21'b111111111111111111110;
		14'b01101111100110:	sigmoid = 21'b111111111111111111110;
		14'b01101111100111:	sigmoid = 21'b111111111111111111110;
		14'b01101111101000:	sigmoid = 21'b111111111111111111110;
		14'b01101111101001:	sigmoid = 21'b111111111111111111110;
		14'b01101111101010:	sigmoid = 21'b111111111111111111110;
		14'b01101111101011:	sigmoid = 21'b111111111111111111110;
		14'b01101111101100:	sigmoid = 21'b111111111111111111110;
		14'b01101111101101:	sigmoid = 21'b111111111111111111110;
		14'b01101111101110:	sigmoid = 21'b111111111111111111110;
		14'b01101111101111:	sigmoid = 21'b111111111111111111110;
		14'b01101111110000:	sigmoid = 21'b111111111111111111110;
		14'b01101111110001:	sigmoid = 21'b111111111111111111110;
		14'b01101111110010:	sigmoid = 21'b111111111111111111110;
		14'b01101111110011:	sigmoid = 21'b111111111111111111110;
		14'b01101111110100:	sigmoid = 21'b111111111111111111110;
		14'b01101111110101:	sigmoid = 21'b111111111111111111110;
		14'b01101111110110:	sigmoid = 21'b111111111111111111110;
		14'b01101111110111:	sigmoid = 21'b111111111111111111110;
		14'b01101111111000:	sigmoid = 21'b111111111111111111110;
		14'b01101111111001:	sigmoid = 21'b111111111111111111110;
		14'b01101111111010:	sigmoid = 21'b111111111111111111110;
		14'b01101111111011:	sigmoid = 21'b111111111111111111110;
		14'b01101111111100:	sigmoid = 21'b111111111111111111110;
		14'b01101111111101:	sigmoid = 21'b111111111111111111110;
		14'b01101111111110:	sigmoid = 21'b111111111111111111110;
		14'b01101111111111:	sigmoid = 21'b111111111111111111110;
		14'b01110000000000:	sigmoid = 21'b111111111111111111110;
		14'b01110000000001:	sigmoid = 21'b111111111111111111110;
		14'b01110000000010:	sigmoid = 21'b111111111111111111110;
		14'b01110000000011:	sigmoid = 21'b111111111111111111110;
		14'b01110000000100:	sigmoid = 21'b111111111111111111110;
		14'b01110000000101:	sigmoid = 21'b111111111111111111110;
		14'b01110000000110:	sigmoid = 21'b111111111111111111110;
		14'b01110000000111:	sigmoid = 21'b111111111111111111110;
		14'b01110000001000:	sigmoid = 21'b111111111111111111110;
		14'b01110000001001:	sigmoid = 21'b111111111111111111110;
		14'b01110000001010:	sigmoid = 21'b111111111111111111110;
		14'b01110000001011:	sigmoid = 21'b111111111111111111110;
		14'b01110000001100:	sigmoid = 21'b111111111111111111110;
		14'b01110000001101:	sigmoid = 21'b111111111111111111110;
		14'b01110000001110:	sigmoid = 21'b111111111111111111110;
		14'b01110000001111:	sigmoid = 21'b111111111111111111110;
		14'b01110000010000:	sigmoid = 21'b111111111111111111110;
		14'b01110000010001:	sigmoid = 21'b111111111111111111110;
		14'b01110000010010:	sigmoid = 21'b111111111111111111110;
		14'b01110000010011:	sigmoid = 21'b111111111111111111110;
		14'b01110000010100:	sigmoid = 21'b111111111111111111110;
		14'b01110000010101:	sigmoid = 21'b111111111111111111110;
		14'b01110000010110:	sigmoid = 21'b111111111111111111110;
		14'b01110000010111:	sigmoid = 21'b111111111111111111110;
		14'b01110000011000:	sigmoid = 21'b111111111111111111110;
		14'b01110000011001:	sigmoid = 21'b111111111111111111110;
		14'b01110000011010:	sigmoid = 21'b111111111111111111110;
		14'b01110000011011:	sigmoid = 21'b111111111111111111110;
		14'b01110000011100:	sigmoid = 21'b111111111111111111110;
		14'b01110000011101:	sigmoid = 21'b111111111111111111110;
		14'b01110000011110:	sigmoid = 21'b111111111111111111110;
		14'b01110000011111:	sigmoid = 21'b111111111111111111110;
		14'b01110000100000:	sigmoid = 21'b111111111111111111110;
		14'b01110000100001:	sigmoid = 21'b111111111111111111110;
		14'b01110000100010:	sigmoid = 21'b111111111111111111110;
		14'b01110000100011:	sigmoid = 21'b111111111111111111110;
		14'b01110000100100:	sigmoid = 21'b111111111111111111110;
		14'b01110000100101:	sigmoid = 21'b111111111111111111110;
		14'b01110000100110:	sigmoid = 21'b111111111111111111110;
		14'b01110000100111:	sigmoid = 21'b111111111111111111110;
		14'b01110000101000:	sigmoid = 21'b111111111111111111110;
		14'b01110000101001:	sigmoid = 21'b111111111111111111110;
		14'b01110000101010:	sigmoid = 21'b111111111111111111110;
		14'b01110000101011:	sigmoid = 21'b111111111111111111110;
		14'b01110000101100:	sigmoid = 21'b111111111111111111110;
		14'b01110000101101:	sigmoid = 21'b111111111111111111110;
		14'b01110000101110:	sigmoid = 21'b111111111111111111110;
		14'b01110000101111:	sigmoid = 21'b111111111111111111110;
		14'b01110000110000:	sigmoid = 21'b111111111111111111110;
		14'b01110000110001:	sigmoid = 21'b111111111111111111110;
		14'b01110000110010:	sigmoid = 21'b111111111111111111110;
		14'b01110000110011:	sigmoid = 21'b111111111111111111110;
		14'b01110000110100:	sigmoid = 21'b111111111111111111110;
		14'b01110000110101:	sigmoid = 21'b111111111111111111110;
		14'b01110000110110:	sigmoid = 21'b111111111111111111110;
		14'b01110000110111:	sigmoid = 21'b111111111111111111110;
		14'b01110000111000:	sigmoid = 21'b111111111111111111110;
		14'b01110000111001:	sigmoid = 21'b111111111111111111110;
		14'b01110000111010:	sigmoid = 21'b111111111111111111110;
		14'b01110000111011:	sigmoid = 21'b111111111111111111110;
		14'b01110000111100:	sigmoid = 21'b111111111111111111110;
		14'b01110000111101:	sigmoid = 21'b111111111111111111110;
		14'b01110000111110:	sigmoid = 21'b111111111111111111110;
		14'b01110000111111:	sigmoid = 21'b111111111111111111110;
		14'b01110001000000:	sigmoid = 21'b111111111111111111110;
		14'b01110001000001:	sigmoid = 21'b111111111111111111110;
		14'b01110001000010:	sigmoid = 21'b111111111111111111110;
		14'b01110001000011:	sigmoid = 21'b111111111111111111110;
		14'b01110001000100:	sigmoid = 21'b111111111111111111110;
		14'b01110001000101:	sigmoid = 21'b111111111111111111110;
		14'b01110001000110:	sigmoid = 21'b111111111111111111110;
		14'b01110001000111:	sigmoid = 21'b111111111111111111110;
		14'b01110001001000:	sigmoid = 21'b111111111111111111110;
		14'b01110001001001:	sigmoid = 21'b111111111111111111110;
		14'b01110001001010:	sigmoid = 21'b111111111111111111110;
		14'b01110001001011:	sigmoid = 21'b111111111111111111110;
		14'b01110001001100:	sigmoid = 21'b111111111111111111110;
		14'b01110001001101:	sigmoid = 21'b111111111111111111110;
		14'b01110001001110:	sigmoid = 21'b111111111111111111110;
		14'b01110001001111:	sigmoid = 21'b111111111111111111110;
		14'b01110001010000:	sigmoid = 21'b111111111111111111110;
		14'b01110001010001:	sigmoid = 21'b111111111111111111110;
		14'b01110001010010:	sigmoid = 21'b111111111111111111110;
		14'b01110001010011:	sigmoid = 21'b111111111111111111110;
		14'b01110001010100:	sigmoid = 21'b111111111111111111110;
		14'b01110001010101:	sigmoid = 21'b111111111111111111110;
		14'b01110001010110:	sigmoid = 21'b111111111111111111110;
		14'b01110001010111:	sigmoid = 21'b111111111111111111110;
		14'b01110001011000:	sigmoid = 21'b111111111111111111110;
		14'b01110001011001:	sigmoid = 21'b111111111111111111110;
		14'b01110001011010:	sigmoid = 21'b111111111111111111110;
		14'b01110001011011:	sigmoid = 21'b111111111111111111110;
		14'b01110001011100:	sigmoid = 21'b111111111111111111110;
		14'b01110001011101:	sigmoid = 21'b111111111111111111110;
		14'b01110001011110:	sigmoid = 21'b111111111111111111110;
		14'b01110001011111:	sigmoid = 21'b111111111111111111110;
		14'b01110001100000:	sigmoid = 21'b111111111111111111110;
		14'b01110001100001:	sigmoid = 21'b111111111111111111110;
		14'b01110001100010:	sigmoid = 21'b111111111111111111110;
		14'b01110001100011:	sigmoid = 21'b111111111111111111110;
		14'b01110001100100:	sigmoid = 21'b111111111111111111110;
		14'b01110001100101:	sigmoid = 21'b111111111111111111110;
		14'b01110001100110:	sigmoid = 21'b111111111111111111110;
		14'b01110001100111:	sigmoid = 21'b111111111111111111110;
		14'b01110001101000:	sigmoid = 21'b111111111111111111110;
		14'b01110001101001:	sigmoid = 21'b111111111111111111110;
		14'b01110001101010:	sigmoid = 21'b111111111111111111110;
		14'b01110001101011:	sigmoid = 21'b111111111111111111110;
		14'b01110001101100:	sigmoid = 21'b111111111111111111110;
		14'b01110001101101:	sigmoid = 21'b111111111111111111110;
		14'b01110001101110:	sigmoid = 21'b111111111111111111110;
		14'b01110001101111:	sigmoid = 21'b111111111111111111110;
		14'b01110001110000:	sigmoid = 21'b111111111111111111110;
		14'b01110001110001:	sigmoid = 21'b111111111111111111110;
		14'b01110001110010:	sigmoid = 21'b111111111111111111110;
		14'b01110001110011:	sigmoid = 21'b111111111111111111110;
		14'b01110001110100:	sigmoid = 21'b111111111111111111110;
		14'b01110001110101:	sigmoid = 21'b111111111111111111110;
		14'b01110001110110:	sigmoid = 21'b111111111111111111110;
		14'b01110001110111:	sigmoid = 21'b111111111111111111110;
		14'b01110001111000:	sigmoid = 21'b111111111111111111110;
		14'b01110001111001:	sigmoid = 21'b111111111111111111110;
		14'b01110001111010:	sigmoid = 21'b111111111111111111110;
		14'b01110001111011:	sigmoid = 21'b111111111111111111110;
		14'b01110001111100:	sigmoid = 21'b111111111111111111110;
		14'b01110001111101:	sigmoid = 21'b111111111111111111110;
		14'b01110001111110:	sigmoid = 21'b111111111111111111110;
		14'b01110001111111:	sigmoid = 21'b111111111111111111110;
		14'b01110010000000:	sigmoid = 21'b111111111111111111110;
		14'b01110010000001:	sigmoid = 21'b111111111111111111110;
		14'b01110010000010:	sigmoid = 21'b111111111111111111110;
		14'b01110010000011:	sigmoid = 21'b111111111111111111110;
		14'b01110010000100:	sigmoid = 21'b111111111111111111110;
		14'b01110010000101:	sigmoid = 21'b111111111111111111110;
		14'b01110010000110:	sigmoid = 21'b111111111111111111110;
		14'b01110010000111:	sigmoid = 21'b111111111111111111110;
		14'b01110010001000:	sigmoid = 21'b111111111111111111110;
		14'b01110010001001:	sigmoid = 21'b111111111111111111110;
		14'b01110010001010:	sigmoid = 21'b111111111111111111110;
		14'b01110010001011:	sigmoid = 21'b111111111111111111110;
		14'b01110010001100:	sigmoid = 21'b111111111111111111110;
		14'b01110010001101:	sigmoid = 21'b111111111111111111110;
		14'b01110010001110:	sigmoid = 21'b111111111111111111110;
		14'b01110010001111:	sigmoid = 21'b111111111111111111110;
		14'b01110010010000:	sigmoid = 21'b111111111111111111110;
		14'b01110010010001:	sigmoid = 21'b111111111111111111110;
		14'b01110010010010:	sigmoid = 21'b111111111111111111110;
		14'b01110010010011:	sigmoid = 21'b111111111111111111110;
		14'b01110010010100:	sigmoid = 21'b111111111111111111110;
		14'b01110010010101:	sigmoid = 21'b111111111111111111110;
		14'b01110010010110:	sigmoid = 21'b111111111111111111110;
		14'b01110010010111:	sigmoid = 21'b111111111111111111110;
		14'b01110010011000:	sigmoid = 21'b111111111111111111110;
		14'b01110010011001:	sigmoid = 21'b111111111111111111110;
		14'b01110010011010:	sigmoid = 21'b111111111111111111110;
		14'b01110010011011:	sigmoid = 21'b111111111111111111110;
		14'b01110010011100:	sigmoid = 21'b111111111111111111110;
		14'b01110010011101:	sigmoid = 21'b111111111111111111110;
		14'b01110010011110:	sigmoid = 21'b111111111111111111110;
		14'b01110010011111:	sigmoid = 21'b111111111111111111110;
		14'b01110010100000:	sigmoid = 21'b111111111111111111110;
		14'b01110010100001:	sigmoid = 21'b111111111111111111110;
		14'b01110010100010:	sigmoid = 21'b111111111111111111110;
		14'b01110010100011:	sigmoid = 21'b111111111111111111110;
		14'b01110010100100:	sigmoid = 21'b111111111111111111110;
		14'b01110010100101:	sigmoid = 21'b111111111111111111110;
		14'b01110010100110:	sigmoid = 21'b111111111111111111110;
		14'b01110010100111:	sigmoid = 21'b111111111111111111110;
		14'b01110010101000:	sigmoid = 21'b111111111111111111110;
		14'b01110010101001:	sigmoid = 21'b111111111111111111110;
		14'b01110010101010:	sigmoid = 21'b111111111111111111110;
		14'b01110010101011:	sigmoid = 21'b111111111111111111110;
		14'b01110010101100:	sigmoid = 21'b111111111111111111110;
		14'b01110010101101:	sigmoid = 21'b111111111111111111110;
		14'b01110010101110:	sigmoid = 21'b111111111111111111110;
		14'b01110010101111:	sigmoid = 21'b111111111111111111110;
		14'b01110010110000:	sigmoid = 21'b111111111111111111110;
		14'b01110010110001:	sigmoid = 21'b111111111111111111110;
		14'b01110010110010:	sigmoid = 21'b111111111111111111110;
		14'b01110010110011:	sigmoid = 21'b111111111111111111110;
		14'b01110010110100:	sigmoid = 21'b111111111111111111110;
		14'b01110010110101:	sigmoid = 21'b111111111111111111110;
		14'b01110010110110:	sigmoid = 21'b111111111111111111110;
		14'b01110010110111:	sigmoid = 21'b111111111111111111110;
		14'b01110010111000:	sigmoid = 21'b111111111111111111110;
		14'b01110010111001:	sigmoid = 21'b111111111111111111110;
		14'b01110010111010:	sigmoid = 21'b111111111111111111110;
		14'b01110010111011:	sigmoid = 21'b111111111111111111110;
		14'b01110010111100:	sigmoid = 21'b111111111111111111110;
		14'b01110010111101:	sigmoid = 21'b111111111111111111110;
		14'b01110010111110:	sigmoid = 21'b111111111111111111110;
		14'b01110010111111:	sigmoid = 21'b111111111111111111110;
		14'b01110011000000:	sigmoid = 21'b111111111111111111110;
		14'b01110011000001:	sigmoid = 21'b111111111111111111110;
		14'b01110011000010:	sigmoid = 21'b111111111111111111110;
		14'b01110011000011:	sigmoid = 21'b111111111111111111110;
		14'b01110011000100:	sigmoid = 21'b111111111111111111110;
		14'b01110011000101:	sigmoid = 21'b111111111111111111110;
		14'b01110011000110:	sigmoid = 21'b111111111111111111110;
		14'b01110011000111:	sigmoid = 21'b111111111111111111110;
		14'b01110011001000:	sigmoid = 21'b111111111111111111110;
		14'b01110011001001:	sigmoid = 21'b111111111111111111110;
		14'b01110011001010:	sigmoid = 21'b111111111111111111110;
		14'b01110011001011:	sigmoid = 21'b111111111111111111110;
		14'b01110011001100:	sigmoid = 21'b111111111111111111110;
		14'b01110011001101:	sigmoid = 21'b111111111111111111110;
		14'b01110011001110:	sigmoid = 21'b111111111111111111110;
		14'b01110011001111:	sigmoid = 21'b111111111111111111110;
		14'b01110011010000:	sigmoid = 21'b111111111111111111110;
		14'b01110011010001:	sigmoid = 21'b111111111111111111110;
		14'b01110011010010:	sigmoid = 21'b111111111111111111110;
		14'b01110011010011:	sigmoid = 21'b111111111111111111110;
		14'b01110011010100:	sigmoid = 21'b111111111111111111110;
		14'b01110011010101:	sigmoid = 21'b111111111111111111110;
		14'b01110011010110:	sigmoid = 21'b111111111111111111110;
		14'b01110011010111:	sigmoid = 21'b111111111111111111110;
		14'b01110011011000:	sigmoid = 21'b111111111111111111110;
		14'b01110011011001:	sigmoid = 21'b111111111111111111110;
		14'b01110011011010:	sigmoid = 21'b111111111111111111110;
		14'b01110011011011:	sigmoid = 21'b111111111111111111110;
		14'b01110011011100:	sigmoid = 21'b111111111111111111110;
		14'b01110011011101:	sigmoid = 21'b111111111111111111110;
		14'b01110011011110:	sigmoid = 21'b111111111111111111110;
		14'b01110011011111:	sigmoid = 21'b111111111111111111110;
		14'b01110011100000:	sigmoid = 21'b111111111111111111110;
		14'b01110011100001:	sigmoid = 21'b111111111111111111110;
		14'b01110011100010:	sigmoid = 21'b111111111111111111110;
		14'b01110011100011:	sigmoid = 21'b111111111111111111110;
		14'b01110011100100:	sigmoid = 21'b111111111111111111110;
		14'b01110011100101:	sigmoid = 21'b111111111111111111110;
		14'b01110011100110:	sigmoid = 21'b111111111111111111110;
		14'b01110011100111:	sigmoid = 21'b111111111111111111110;
		14'b01110011101000:	sigmoid = 21'b111111111111111111110;
		14'b01110011101001:	sigmoid = 21'b111111111111111111110;
		14'b01110011101010:	sigmoid = 21'b111111111111111111110;
		14'b01110011101011:	sigmoid = 21'b111111111111111111110;
		14'b01110011101100:	sigmoid = 21'b111111111111111111110;
		14'b01110011101101:	sigmoid = 21'b111111111111111111110;
		14'b01110011101110:	sigmoid = 21'b111111111111111111110;
		14'b01110011101111:	sigmoid = 21'b111111111111111111110;
		14'b01110011110000:	sigmoid = 21'b111111111111111111110;
		14'b01110011110001:	sigmoid = 21'b111111111111111111110;
		14'b01110011110010:	sigmoid = 21'b111111111111111111110;
		14'b01110011110011:	sigmoid = 21'b111111111111111111110;
		14'b01110011110100:	sigmoid = 21'b111111111111111111110;
		14'b01110011110101:	sigmoid = 21'b111111111111111111110;
		14'b01110011110110:	sigmoid = 21'b111111111111111111110;
		14'b01110011110111:	sigmoid = 21'b111111111111111111110;
		14'b01110011111000:	sigmoid = 21'b111111111111111111110;
		14'b01110011111001:	sigmoid = 21'b111111111111111111110;
		14'b01110011111010:	sigmoid = 21'b111111111111111111110;
		14'b01110011111011:	sigmoid = 21'b111111111111111111110;
		14'b01110011111100:	sigmoid = 21'b111111111111111111110;
		14'b01110011111101:	sigmoid = 21'b111111111111111111110;
		14'b01110011111110:	sigmoid = 21'b111111111111111111110;
		14'b01110011111111:	sigmoid = 21'b111111111111111111110;
		14'b01110100000000:	sigmoid = 21'b111111111111111111110;
		14'b01110100000001:	sigmoid = 21'b111111111111111111110;
		14'b01110100000010:	sigmoid = 21'b111111111111111111110;
		14'b01110100000011:	sigmoid = 21'b111111111111111111110;
		14'b01110100000100:	sigmoid = 21'b111111111111111111110;
		14'b01110100000101:	sigmoid = 21'b111111111111111111110;
		14'b01110100000110:	sigmoid = 21'b111111111111111111110;
		14'b01110100000111:	sigmoid = 21'b111111111111111111110;
		14'b01110100001000:	sigmoid = 21'b111111111111111111110;
		14'b01110100001001:	sigmoid = 21'b111111111111111111110;
		14'b01110100001010:	sigmoid = 21'b111111111111111111110;
		14'b01110100001011:	sigmoid = 21'b111111111111111111110;
		14'b01110100001100:	sigmoid = 21'b111111111111111111110;
		14'b01110100001101:	sigmoid = 21'b111111111111111111110;
		14'b01110100001110:	sigmoid = 21'b111111111111111111110;
		14'b01110100001111:	sigmoid = 21'b111111111111111111110;
		14'b01110100010000:	sigmoid = 21'b111111111111111111110;
		14'b01110100010001:	sigmoid = 21'b111111111111111111110;
		14'b01110100010010:	sigmoid = 21'b111111111111111111110;
		14'b01110100010011:	sigmoid = 21'b111111111111111111110;
		14'b01110100010100:	sigmoid = 21'b111111111111111111110;
		14'b01110100010101:	sigmoid = 21'b111111111111111111110;
		14'b01110100010110:	sigmoid = 21'b111111111111111111110;
		14'b01110100010111:	sigmoid = 21'b111111111111111111110;
		14'b01110100011000:	sigmoid = 21'b111111111111111111110;
		14'b01110100011001:	sigmoid = 21'b111111111111111111110;
		14'b01110100011010:	sigmoid = 21'b111111111111111111110;
		14'b01110100011011:	sigmoid = 21'b111111111111111111110;
		14'b01110100011100:	sigmoid = 21'b111111111111111111110;
		14'b01110100011101:	sigmoid = 21'b111111111111111111111;
		14'b01110100011110:	sigmoid = 21'b111111111111111111111;
		14'b01110100011111:	sigmoid = 21'b111111111111111111111;
		14'b01110100100000:	sigmoid = 21'b111111111111111111111;
		14'b01110100100001:	sigmoid = 21'b111111111111111111111;
		14'b01110100100010:	sigmoid = 21'b111111111111111111111;
		14'b01110100100011:	sigmoid = 21'b111111111111111111111;
		14'b01110100100100:	sigmoid = 21'b111111111111111111111;
		14'b01110100100101:	sigmoid = 21'b111111111111111111111;
		14'b01110100100110:	sigmoid = 21'b111111111111111111111;
		14'b01110100100111:	sigmoid = 21'b111111111111111111111;
		14'b01110100101000:	sigmoid = 21'b111111111111111111111;
		14'b01110100101001:	sigmoid = 21'b111111111111111111111;
		14'b01110100101010:	sigmoid = 21'b111111111111111111111;
		14'b01110100101011:	sigmoid = 21'b111111111111111111111;
		14'b01110100101100:	sigmoid = 21'b111111111111111111111;
		14'b01110100101101:	sigmoid = 21'b111111111111111111111;
		14'b01110100101110:	sigmoid = 21'b111111111111111111111;
		14'b01110100101111:	sigmoid = 21'b111111111111111111111;
		14'b01110100110000:	sigmoid = 21'b111111111111111111111;
		14'b01110100110001:	sigmoid = 21'b111111111111111111111;
		14'b01110100110010:	sigmoid = 21'b111111111111111111111;
		14'b01110100110011:	sigmoid = 21'b111111111111111111111;
		14'b01110100110100:	sigmoid = 21'b111111111111111111111;
		14'b01110100110101:	sigmoid = 21'b111111111111111111111;
		14'b01110100110110:	sigmoid = 21'b111111111111111111111;
		14'b01110100110111:	sigmoid = 21'b111111111111111111111;
		14'b01110100111000:	sigmoid = 21'b111111111111111111111;
		14'b01110100111001:	sigmoid = 21'b111111111111111111111;
		14'b01110100111010:	sigmoid = 21'b111111111111111111111;
		14'b01110100111011:	sigmoid = 21'b111111111111111111111;
		14'b01110100111100:	sigmoid = 21'b111111111111111111111;
		14'b01110100111101:	sigmoid = 21'b111111111111111111111;
		14'b01110100111110:	sigmoid = 21'b111111111111111111111;
		14'b01110100111111:	sigmoid = 21'b111111111111111111111;
		14'b01110101000000:	sigmoid = 21'b111111111111111111111;
		14'b01110101000001:	sigmoid = 21'b111111111111111111111;
		14'b01110101000010:	sigmoid = 21'b111111111111111111111;
		14'b01110101000011:	sigmoid = 21'b111111111111111111111;
		14'b01110101000100:	sigmoid = 21'b111111111111111111111;
		14'b01110101000101:	sigmoid = 21'b111111111111111111111;
		14'b01110101000110:	sigmoid = 21'b111111111111111111111;
		14'b01110101000111:	sigmoid = 21'b111111111111111111111;
		14'b01110101001000:	sigmoid = 21'b111111111111111111111;
		14'b01110101001001:	sigmoid = 21'b111111111111111111111;
		14'b01110101001010:	sigmoid = 21'b111111111111111111111;
		14'b01110101001011:	sigmoid = 21'b111111111111111111111;
		14'b01110101001100:	sigmoid = 21'b111111111111111111111;
		14'b01110101001101:	sigmoid = 21'b111111111111111111111;
		14'b01110101001110:	sigmoid = 21'b111111111111111111111;
		14'b01110101001111:	sigmoid = 21'b111111111111111111111;
		14'b01110101010000:	sigmoid = 21'b111111111111111111111;
		14'b01110101010001:	sigmoid = 21'b111111111111111111111;
		14'b01110101010010:	sigmoid = 21'b111111111111111111111;
		14'b01110101010011:	sigmoid = 21'b111111111111111111111;
		14'b01110101010100:	sigmoid = 21'b111111111111111111111;
		14'b01110101010101:	sigmoid = 21'b111111111111111111111;
		14'b01110101010110:	sigmoid = 21'b111111111111111111111;
		14'b01110101010111:	sigmoid = 21'b111111111111111111111;
		14'b01110101011000:	sigmoid = 21'b111111111111111111111;
		14'b01110101011001:	sigmoid = 21'b111111111111111111111;
		14'b01110101011010:	sigmoid = 21'b111111111111111111111;
		14'b01110101011011:	sigmoid = 21'b111111111111111111111;
		14'b01110101011100:	sigmoid = 21'b111111111111111111111;
		14'b01110101011101:	sigmoid = 21'b111111111111111111111;
		14'b01110101011110:	sigmoid = 21'b111111111111111111111;
		14'b01110101011111:	sigmoid = 21'b111111111111111111111;
		14'b01110101100000:	sigmoid = 21'b111111111111111111111;
		14'b01110101100001:	sigmoid = 21'b111111111111111111111;
		14'b01110101100010:	sigmoid = 21'b111111111111111111111;
		14'b01110101100011:	sigmoid = 21'b111111111111111111111;
		14'b01110101100100:	sigmoid = 21'b111111111111111111111;
		14'b01110101100101:	sigmoid = 21'b111111111111111111111;
		14'b01110101100110:	sigmoid = 21'b111111111111111111111;
		14'b01110101100111:	sigmoid = 21'b111111111111111111111;
		14'b01110101101000:	sigmoid = 21'b111111111111111111111;
		14'b01110101101001:	sigmoid = 21'b111111111111111111111;
		14'b01110101101010:	sigmoid = 21'b111111111111111111111;
		14'b01110101101011:	sigmoid = 21'b111111111111111111111;
		14'b01110101101100:	sigmoid = 21'b111111111111111111111;
		14'b01110101101101:	sigmoid = 21'b111111111111111111111;
		14'b01110101101110:	sigmoid = 21'b111111111111111111111;
		14'b01110101101111:	sigmoid = 21'b111111111111111111111;
		14'b01110101110000:	sigmoid = 21'b111111111111111111111;
		14'b01110101110001:	sigmoid = 21'b111111111111111111111;
		14'b01110101110010:	sigmoid = 21'b111111111111111111111;
		14'b01110101110011:	sigmoid = 21'b111111111111111111111;
		14'b01110101110100:	sigmoid = 21'b111111111111111111111;
		14'b01110101110101:	sigmoid = 21'b111111111111111111111;
		14'b01110101110110:	sigmoid = 21'b111111111111111111111;
		14'b01110101110111:	sigmoid = 21'b111111111111111111111;
		14'b01110101111000:	sigmoid = 21'b111111111111111111111;
		14'b01110101111001:	sigmoid = 21'b111111111111111111111;
		14'b01110101111010:	sigmoid = 21'b111111111111111111111;
		14'b01110101111011:	sigmoid = 21'b111111111111111111111;
		14'b01110101111100:	sigmoid = 21'b111111111111111111111;
		14'b01110101111101:	sigmoid = 21'b111111111111111111111;
		14'b01110101111110:	sigmoid = 21'b111111111111111111111;
		14'b01110101111111:	sigmoid = 21'b111111111111111111111;
		14'b01110110000000:	sigmoid = 21'b111111111111111111111;
		14'b01110110000001:	sigmoid = 21'b111111111111111111111;
		14'b01110110000010:	sigmoid = 21'b111111111111111111111;
		14'b01110110000011:	sigmoid = 21'b111111111111111111111;
		14'b01110110000100:	sigmoid = 21'b111111111111111111111;
		14'b01110110000101:	sigmoid = 21'b111111111111111111111;
		14'b01110110000110:	sigmoid = 21'b111111111111111111111;
		14'b01110110000111:	sigmoid = 21'b111111111111111111111;
		14'b01110110001000:	sigmoid = 21'b111111111111111111111;
		14'b01110110001001:	sigmoid = 21'b111111111111111111111;
		14'b01110110001010:	sigmoid = 21'b111111111111111111111;
		14'b01110110001011:	sigmoid = 21'b111111111111111111111;
		14'b01110110001100:	sigmoid = 21'b111111111111111111111;
		14'b01110110001101:	sigmoid = 21'b111111111111111111111;
		14'b01110110001110:	sigmoid = 21'b111111111111111111111;
		14'b01110110001111:	sigmoid = 21'b111111111111111111111;
		14'b01110110010000:	sigmoid = 21'b111111111111111111111;
		14'b01110110010001:	sigmoid = 21'b111111111111111111111;
		14'b01110110010010:	sigmoid = 21'b111111111111111111111;
		14'b01110110010011:	sigmoid = 21'b111111111111111111111;
		14'b01110110010100:	sigmoid = 21'b111111111111111111111;
		14'b01110110010101:	sigmoid = 21'b111111111111111111111;
		14'b01110110010110:	sigmoid = 21'b111111111111111111111;
		14'b01110110010111:	sigmoid = 21'b111111111111111111111;
		14'b01110110011000:	sigmoid = 21'b111111111111111111111;
		14'b01110110011001:	sigmoid = 21'b111111111111111111111;
		14'b01110110011010:	sigmoid = 21'b111111111111111111111;
		14'b01110110011011:	sigmoid = 21'b111111111111111111111;
		14'b01110110011100:	sigmoid = 21'b111111111111111111111;
		14'b01110110011101:	sigmoid = 21'b111111111111111111111;
		14'b01110110011110:	sigmoid = 21'b111111111111111111111;
		14'b01110110011111:	sigmoid = 21'b111111111111111111111;
		14'b01110110100000:	sigmoid = 21'b111111111111111111111;
		14'b01110110100001:	sigmoid = 21'b111111111111111111111;
		14'b01110110100010:	sigmoid = 21'b111111111111111111111;
		14'b01110110100011:	sigmoid = 21'b111111111111111111111;
		14'b01110110100100:	sigmoid = 21'b111111111111111111111;
		14'b01110110100101:	sigmoid = 21'b111111111111111111111;
		14'b01110110100110:	sigmoid = 21'b111111111111111111111;
		14'b01110110100111:	sigmoid = 21'b111111111111111111111;
		14'b01110110101000:	sigmoid = 21'b111111111111111111111;
		14'b01110110101001:	sigmoid = 21'b111111111111111111111;
		14'b01110110101010:	sigmoid = 21'b111111111111111111111;
		14'b01110110101011:	sigmoid = 21'b111111111111111111111;
		14'b01110110101100:	sigmoid = 21'b111111111111111111111;
		14'b01110110101101:	sigmoid = 21'b111111111111111111111;
		14'b01110110101110:	sigmoid = 21'b111111111111111111111;
		14'b01110110101111:	sigmoid = 21'b111111111111111111111;
		14'b01110110110000:	sigmoid = 21'b111111111111111111111;
		14'b01110110110001:	sigmoid = 21'b111111111111111111111;
		14'b01110110110010:	sigmoid = 21'b111111111111111111111;
		14'b01110110110011:	sigmoid = 21'b111111111111111111111;
		14'b01110110110100:	sigmoid = 21'b111111111111111111111;
		14'b01110110110101:	sigmoid = 21'b111111111111111111111;
		14'b01110110110110:	sigmoid = 21'b111111111111111111111;
		14'b01110110110111:	sigmoid = 21'b111111111111111111111;
		14'b01110110111000:	sigmoid = 21'b111111111111111111111;
		14'b01110110111001:	sigmoid = 21'b111111111111111111111;
		14'b01110110111010:	sigmoid = 21'b111111111111111111111;
		14'b01110110111011:	sigmoid = 21'b111111111111111111111;
		14'b01110110111100:	sigmoid = 21'b111111111111111111111;
		14'b01110110111101:	sigmoid = 21'b111111111111111111111;
		14'b01110110111110:	sigmoid = 21'b111111111111111111111;
		14'b01110110111111:	sigmoid = 21'b111111111111111111111;
		14'b01110111000000:	sigmoid = 21'b111111111111111111111;
		14'b01110111000001:	sigmoid = 21'b111111111111111111111;
		14'b01110111000010:	sigmoid = 21'b111111111111111111111;
		14'b01110111000011:	sigmoid = 21'b111111111111111111111;
		14'b01110111000100:	sigmoid = 21'b111111111111111111111;
		14'b01110111000101:	sigmoid = 21'b111111111111111111111;
		14'b01110111000110:	sigmoid = 21'b111111111111111111111;
		14'b01110111000111:	sigmoid = 21'b111111111111111111111;
		14'b01110111001000:	sigmoid = 21'b111111111111111111111;
		14'b01110111001001:	sigmoid = 21'b111111111111111111111;
		14'b01110111001010:	sigmoid = 21'b111111111111111111111;
		14'b01110111001011:	sigmoid = 21'b111111111111111111111;
		14'b01110111001100:	sigmoid = 21'b111111111111111111111;
		14'b01110111001101:	sigmoid = 21'b111111111111111111111;
		14'b01110111001110:	sigmoid = 21'b111111111111111111111;
		14'b01110111001111:	sigmoid = 21'b111111111111111111111;
		14'b01110111010000:	sigmoid = 21'b111111111111111111111;
		14'b01110111010001:	sigmoid = 21'b111111111111111111111;
		14'b01110111010010:	sigmoid = 21'b111111111111111111111;
		14'b01110111010011:	sigmoid = 21'b111111111111111111111;
		14'b01110111010100:	sigmoid = 21'b111111111111111111111;
		14'b01110111010101:	sigmoid = 21'b111111111111111111111;
		14'b01110111010110:	sigmoid = 21'b111111111111111111111;
		14'b01110111010111:	sigmoid = 21'b111111111111111111111;
		14'b01110111011000:	sigmoid = 21'b111111111111111111111;
		14'b01110111011001:	sigmoid = 21'b111111111111111111111;
		14'b01110111011010:	sigmoid = 21'b111111111111111111111;
		14'b01110111011011:	sigmoid = 21'b111111111111111111111;
		14'b01110111011100:	sigmoid = 21'b111111111111111111111;
		14'b01110111011101:	sigmoid = 21'b111111111111111111111;
		14'b01110111011110:	sigmoid = 21'b111111111111111111111;
		14'b01110111011111:	sigmoid = 21'b111111111111111111111;
		14'b01110111100000:	sigmoid = 21'b111111111111111111111;
		14'b01110111100001:	sigmoid = 21'b111111111111111111111;
		14'b01110111100010:	sigmoid = 21'b111111111111111111111;
		14'b01110111100011:	sigmoid = 21'b111111111111111111111;
		14'b01110111100100:	sigmoid = 21'b111111111111111111111;
		14'b01110111100101:	sigmoid = 21'b111111111111111111111;
		14'b01110111100110:	sigmoid = 21'b111111111111111111111;
		14'b01110111100111:	sigmoid = 21'b111111111111111111111;
		14'b01110111101000:	sigmoid = 21'b111111111111111111111;
		14'b01110111101001:	sigmoid = 21'b111111111111111111111;
		14'b01110111101010:	sigmoid = 21'b111111111111111111111;
		14'b01110111101011:	sigmoid = 21'b111111111111111111111;
		14'b01110111101100:	sigmoid = 21'b111111111111111111111;
		14'b01110111101101:	sigmoid = 21'b111111111111111111111;
		14'b01110111101110:	sigmoid = 21'b111111111111111111111;
		14'b01110111101111:	sigmoid = 21'b111111111111111111111;
		14'b01110111110000:	sigmoid = 21'b111111111111111111111;
		14'b01110111110001:	sigmoid = 21'b111111111111111111111;
		14'b01110111110010:	sigmoid = 21'b111111111111111111111;
		14'b01110111110011:	sigmoid = 21'b111111111111111111111;
		14'b01110111110100:	sigmoid = 21'b111111111111111111111;
		14'b01110111110101:	sigmoid = 21'b111111111111111111111;
		14'b01110111110110:	sigmoid = 21'b111111111111111111111;
		14'b01110111110111:	sigmoid = 21'b111111111111111111111;
		14'b01110111111000:	sigmoid = 21'b111111111111111111111;
		14'b01110111111001:	sigmoid = 21'b111111111111111111111;
		14'b01110111111010:	sigmoid = 21'b111111111111111111111;
		14'b01110111111011:	sigmoid = 21'b111111111111111111111;
		14'b01110111111100:	sigmoid = 21'b111111111111111111111;
		14'b01110111111101:	sigmoid = 21'b111111111111111111111;
		14'b01110111111110:	sigmoid = 21'b111111111111111111111;
		14'b01110111111111:	sigmoid = 21'b111111111111111111111;
		14'b01111000000000:	sigmoid = 21'b111111111111111111111;
		14'b01111000000001:	sigmoid = 21'b111111111111111111111;
		14'b01111000000010:	sigmoid = 21'b111111111111111111111;
		14'b01111000000011:	sigmoid = 21'b111111111111111111111;
		14'b01111000000100:	sigmoid = 21'b111111111111111111111;
		14'b01111000000101:	sigmoid = 21'b111111111111111111111;
		14'b01111000000110:	sigmoid = 21'b111111111111111111111;
		14'b01111000000111:	sigmoid = 21'b111111111111111111111;
		14'b01111000001000:	sigmoid = 21'b111111111111111111111;
		14'b01111000001001:	sigmoid = 21'b111111111111111111111;
		14'b01111000001010:	sigmoid = 21'b111111111111111111111;
		14'b01111000001011:	sigmoid = 21'b111111111111111111111;
		14'b01111000001100:	sigmoid = 21'b111111111111111111111;
		14'b01111000001101:	sigmoid = 21'b111111111111111111111;
		14'b01111000001110:	sigmoid = 21'b111111111111111111111;
		14'b01111000001111:	sigmoid = 21'b111111111111111111111;
		14'b01111000010000:	sigmoid = 21'b111111111111111111111;
		14'b01111000010001:	sigmoid = 21'b111111111111111111111;
		14'b01111000010010:	sigmoid = 21'b111111111111111111111;
		14'b01111000010011:	sigmoid = 21'b111111111111111111111;
		14'b01111000010100:	sigmoid = 21'b111111111111111111111;
		14'b01111000010101:	sigmoid = 21'b111111111111111111111;
		14'b01111000010110:	sigmoid = 21'b111111111111111111111;
		14'b01111000010111:	sigmoid = 21'b111111111111111111111;
		14'b01111000011000:	sigmoid = 21'b111111111111111111111;
		14'b01111000011001:	sigmoid = 21'b111111111111111111111;
		14'b01111000011010:	sigmoid = 21'b111111111111111111111;
		14'b01111000011011:	sigmoid = 21'b111111111111111111111;
		14'b01111000011100:	sigmoid = 21'b111111111111111111111;
		14'b01111000011101:	sigmoid = 21'b111111111111111111111;
		14'b01111000011110:	sigmoid = 21'b111111111111111111111;
		14'b01111000011111:	sigmoid = 21'b111111111111111111111;
		14'b01111000100000:	sigmoid = 21'b111111111111111111111;
		14'b01111000100001:	sigmoid = 21'b111111111111111111111;
		14'b01111000100010:	sigmoid = 21'b111111111111111111111;
		14'b01111000100011:	sigmoid = 21'b111111111111111111111;
		14'b01111000100100:	sigmoid = 21'b111111111111111111111;
		14'b01111000100101:	sigmoid = 21'b111111111111111111111;
		14'b01111000100110:	sigmoid = 21'b111111111111111111111;
		14'b01111000100111:	sigmoid = 21'b111111111111111111111;
		14'b01111000101000:	sigmoid = 21'b111111111111111111111;
		14'b01111000101001:	sigmoid = 21'b111111111111111111111;
		14'b01111000101010:	sigmoid = 21'b111111111111111111111;
		14'b01111000101011:	sigmoid = 21'b111111111111111111111;
		14'b01111000101100:	sigmoid = 21'b111111111111111111111;
		14'b01111000101101:	sigmoid = 21'b111111111111111111111;
		14'b01111000101110:	sigmoid = 21'b111111111111111111111;
		14'b01111000101111:	sigmoid = 21'b111111111111111111111;
		14'b01111000110000:	sigmoid = 21'b111111111111111111111;
		14'b01111000110001:	sigmoid = 21'b111111111111111111111;
		14'b01111000110010:	sigmoid = 21'b111111111111111111111;
		14'b01111000110011:	sigmoid = 21'b111111111111111111111;
		14'b01111000110100:	sigmoid = 21'b111111111111111111111;
		14'b01111000110101:	sigmoid = 21'b111111111111111111111;
		14'b01111000110110:	sigmoid = 21'b111111111111111111111;
		14'b01111000110111:	sigmoid = 21'b111111111111111111111;
		14'b01111000111000:	sigmoid = 21'b111111111111111111111;
		14'b01111000111001:	sigmoid = 21'b111111111111111111111;
		14'b01111000111010:	sigmoid = 21'b111111111111111111111;
		14'b01111000111011:	sigmoid = 21'b111111111111111111111;
		14'b01111000111100:	sigmoid = 21'b111111111111111111111;
		14'b01111000111101:	sigmoid = 21'b111111111111111111111;
		14'b01111000111110:	sigmoid = 21'b111111111111111111111;
		14'b01111000111111:	sigmoid = 21'b111111111111111111111;
		14'b01111001000000:	sigmoid = 21'b111111111111111111111;
		14'b01111001000001:	sigmoid = 21'b111111111111111111111;
		14'b01111001000010:	sigmoid = 21'b111111111111111111111;
		14'b01111001000011:	sigmoid = 21'b111111111111111111111;
		14'b01111001000100:	sigmoid = 21'b111111111111111111111;
		14'b01111001000101:	sigmoid = 21'b111111111111111111111;
		14'b01111001000110:	sigmoid = 21'b111111111111111111111;
		14'b01111001000111:	sigmoid = 21'b111111111111111111111;
		14'b01111001001000:	sigmoid = 21'b111111111111111111111;
		14'b01111001001001:	sigmoid = 21'b111111111111111111111;
		14'b01111001001010:	sigmoid = 21'b111111111111111111111;
		14'b01111001001011:	sigmoid = 21'b111111111111111111111;
		14'b01111001001100:	sigmoid = 21'b111111111111111111111;
		14'b01111001001101:	sigmoid = 21'b111111111111111111111;
		14'b01111001001110:	sigmoid = 21'b111111111111111111111;
		14'b01111001001111:	sigmoid = 21'b111111111111111111111;
		14'b01111001010000:	sigmoid = 21'b111111111111111111111;
		14'b01111001010001:	sigmoid = 21'b111111111111111111111;
		14'b01111001010010:	sigmoid = 21'b111111111111111111111;
		14'b01111001010011:	sigmoid = 21'b111111111111111111111;
		14'b01111001010100:	sigmoid = 21'b111111111111111111111;
		14'b01111001010101:	sigmoid = 21'b111111111111111111111;
		14'b01111001010110:	sigmoid = 21'b111111111111111111111;
		14'b01111001010111:	sigmoid = 21'b111111111111111111111;
		14'b01111001011000:	sigmoid = 21'b111111111111111111111;
		14'b01111001011001:	sigmoid = 21'b111111111111111111111;
		14'b01111001011010:	sigmoid = 21'b111111111111111111111;
		14'b01111001011011:	sigmoid = 21'b111111111111111111111;
		14'b01111001011100:	sigmoid = 21'b111111111111111111111;
		14'b01111001011101:	sigmoid = 21'b111111111111111111111;
		14'b01111001011110:	sigmoid = 21'b111111111111111111111;
		14'b01111001011111:	sigmoid = 21'b111111111111111111111;
		14'b01111001100000:	sigmoid = 21'b111111111111111111111;
		14'b01111001100001:	sigmoid = 21'b111111111111111111111;
		14'b01111001100010:	sigmoid = 21'b111111111111111111111;
		14'b01111001100011:	sigmoid = 21'b111111111111111111111;
		14'b01111001100100:	sigmoid = 21'b111111111111111111111;
		14'b01111001100101:	sigmoid = 21'b111111111111111111111;
		14'b01111001100110:	sigmoid = 21'b111111111111111111111;
		14'b01111001100111:	sigmoid = 21'b111111111111111111111;
		14'b01111001101000:	sigmoid = 21'b111111111111111111111;
		14'b01111001101001:	sigmoid = 21'b111111111111111111111;
		14'b01111001101010:	sigmoid = 21'b111111111111111111111;
		14'b01111001101011:	sigmoid = 21'b111111111111111111111;
		14'b01111001101100:	sigmoid = 21'b111111111111111111111;
		14'b01111001101101:	sigmoid = 21'b111111111111111111111;
		14'b01111001101110:	sigmoid = 21'b111111111111111111111;
		14'b01111001101111:	sigmoid = 21'b111111111111111111111;
		14'b01111001110000:	sigmoid = 21'b111111111111111111111;
		14'b01111001110001:	sigmoid = 21'b111111111111111111111;
		14'b01111001110010:	sigmoid = 21'b111111111111111111111;
		14'b01111001110011:	sigmoid = 21'b111111111111111111111;
		14'b01111001110100:	sigmoid = 21'b111111111111111111111;
		14'b01111001110101:	sigmoid = 21'b111111111111111111111;
		14'b01111001110110:	sigmoid = 21'b111111111111111111111;
		14'b01111001110111:	sigmoid = 21'b111111111111111111111;
		14'b01111001111000:	sigmoid = 21'b111111111111111111111;
		14'b01111001111001:	sigmoid = 21'b111111111111111111111;
		14'b01111001111010:	sigmoid = 21'b111111111111111111111;
		14'b01111001111011:	sigmoid = 21'b111111111111111111111;
		14'b01111001111100:	sigmoid = 21'b111111111111111111111;
		14'b01111001111101:	sigmoid = 21'b111111111111111111111;
		14'b01111001111110:	sigmoid = 21'b111111111111111111111;
		14'b01111001111111:	sigmoid = 21'b111111111111111111111;
		14'b01111010000000:	sigmoid = 21'b111111111111111111111;
		14'b01111010000001:	sigmoid = 21'b111111111111111111111;
		14'b01111010000010:	sigmoid = 21'b111111111111111111111;
		14'b01111010000011:	sigmoid = 21'b111111111111111111111;
		14'b01111010000100:	sigmoid = 21'b111111111111111111111;
		14'b01111010000101:	sigmoid = 21'b111111111111111111111;
		14'b01111010000110:	sigmoid = 21'b111111111111111111111;
		14'b01111010000111:	sigmoid = 21'b111111111111111111111;
		14'b01111010001000:	sigmoid = 21'b111111111111111111111;
		14'b01111010001001:	sigmoid = 21'b111111111111111111111;
		14'b01111010001010:	sigmoid = 21'b111111111111111111111;
		14'b01111010001011:	sigmoid = 21'b111111111111111111111;
		14'b01111010001100:	sigmoid = 21'b111111111111111111111;
		14'b01111010001101:	sigmoid = 21'b111111111111111111111;
		14'b01111010001110:	sigmoid = 21'b111111111111111111111;
		14'b01111010001111:	sigmoid = 21'b111111111111111111111;
		14'b01111010010000:	sigmoid = 21'b111111111111111111111;
		14'b01111010010001:	sigmoid = 21'b111111111111111111111;
		14'b01111010010010:	sigmoid = 21'b111111111111111111111;
		14'b01111010010011:	sigmoid = 21'b111111111111111111111;
		14'b01111010010100:	sigmoid = 21'b111111111111111111111;
		14'b01111010010101:	sigmoid = 21'b111111111111111111111;
		14'b01111010010110:	sigmoid = 21'b111111111111111111111;
		14'b01111010010111:	sigmoid = 21'b111111111111111111111;
		14'b01111010011000:	sigmoid = 21'b111111111111111111111;
		14'b01111010011001:	sigmoid = 21'b111111111111111111111;
		14'b01111010011010:	sigmoid = 21'b111111111111111111111;
		14'b01111010011011:	sigmoid = 21'b111111111111111111111;
		14'b01111010011100:	sigmoid = 21'b111111111111111111111;
		14'b01111010011101:	sigmoid = 21'b111111111111111111111;
		14'b01111010011110:	sigmoid = 21'b111111111111111111111;
		14'b01111010011111:	sigmoid = 21'b111111111111111111111;
		14'b01111010100000:	sigmoid = 21'b111111111111111111111;
		14'b01111010100001:	sigmoid = 21'b111111111111111111111;
		14'b01111010100010:	sigmoid = 21'b111111111111111111111;
		14'b01111010100011:	sigmoid = 21'b111111111111111111111;
		14'b01111010100100:	sigmoid = 21'b111111111111111111111;
		14'b01111010100101:	sigmoid = 21'b111111111111111111111;
		14'b01111010100110:	sigmoid = 21'b111111111111111111111;
		14'b01111010100111:	sigmoid = 21'b111111111111111111111;
		14'b01111010101000:	sigmoid = 21'b111111111111111111111;
		14'b01111010101001:	sigmoid = 21'b111111111111111111111;
		14'b01111010101010:	sigmoid = 21'b111111111111111111111;
		14'b01111010101011:	sigmoid = 21'b111111111111111111111;
		14'b01111010101100:	sigmoid = 21'b111111111111111111111;
		14'b01111010101101:	sigmoid = 21'b111111111111111111111;
		14'b01111010101110:	sigmoid = 21'b111111111111111111111;
		14'b01111010101111:	sigmoid = 21'b111111111111111111111;
		14'b01111010110000:	sigmoid = 21'b111111111111111111111;
		14'b01111010110001:	sigmoid = 21'b111111111111111111111;
		14'b01111010110010:	sigmoid = 21'b111111111111111111111;
		14'b01111010110011:	sigmoid = 21'b111111111111111111111;
		14'b01111010110100:	sigmoid = 21'b111111111111111111111;
		14'b01111010110101:	sigmoid = 21'b111111111111111111111;
		14'b01111010110110:	sigmoid = 21'b111111111111111111111;
		14'b01111010110111:	sigmoid = 21'b111111111111111111111;
		14'b01111010111000:	sigmoid = 21'b111111111111111111111;
		14'b01111010111001:	sigmoid = 21'b111111111111111111111;
		14'b01111010111010:	sigmoid = 21'b111111111111111111111;
		14'b01111010111011:	sigmoid = 21'b111111111111111111111;
		14'b01111010111100:	sigmoid = 21'b111111111111111111111;
		14'b01111010111101:	sigmoid = 21'b111111111111111111111;
		14'b01111010111110:	sigmoid = 21'b111111111111111111111;
		14'b01111010111111:	sigmoid = 21'b111111111111111111111;
		14'b01111011000000:	sigmoid = 21'b111111111111111111111;
		14'b01111011000001:	sigmoid = 21'b111111111111111111111;
		14'b01111011000010:	sigmoid = 21'b111111111111111111111;
		14'b01111011000011:	sigmoid = 21'b111111111111111111111;
		14'b01111011000100:	sigmoid = 21'b111111111111111111111;
		14'b01111011000101:	sigmoid = 21'b111111111111111111111;
		14'b01111011000110:	sigmoid = 21'b111111111111111111111;
		14'b01111011000111:	sigmoid = 21'b111111111111111111111;
		14'b01111011001000:	sigmoid = 21'b111111111111111111111;
		14'b01111011001001:	sigmoid = 21'b111111111111111111111;
		14'b01111011001010:	sigmoid = 21'b111111111111111111111;
		14'b01111011001011:	sigmoid = 21'b111111111111111111111;
		14'b01111011001100:	sigmoid = 21'b111111111111111111111;
		14'b01111011001101:	sigmoid = 21'b111111111111111111111;
		14'b01111011001110:	sigmoid = 21'b111111111111111111111;
		14'b01111011001111:	sigmoid = 21'b111111111111111111111;
		14'b01111011010000:	sigmoid = 21'b111111111111111111111;
		14'b01111011010001:	sigmoid = 21'b111111111111111111111;
		14'b01111011010010:	sigmoid = 21'b111111111111111111111;
		14'b01111011010011:	sigmoid = 21'b111111111111111111111;
		14'b01111011010100:	sigmoid = 21'b111111111111111111111;
		14'b01111011010101:	sigmoid = 21'b111111111111111111111;
		14'b01111011010110:	sigmoid = 21'b111111111111111111111;
		14'b01111011010111:	sigmoid = 21'b111111111111111111111;
		14'b01111011011000:	sigmoid = 21'b111111111111111111111;
		14'b01111011011001:	sigmoid = 21'b111111111111111111111;
		14'b01111011011010:	sigmoid = 21'b111111111111111111111;
		14'b01111011011011:	sigmoid = 21'b111111111111111111111;
		14'b01111011011100:	sigmoid = 21'b111111111111111111111;
		14'b01111011011101:	sigmoid = 21'b111111111111111111111;
		14'b01111011011110:	sigmoid = 21'b111111111111111111111;
		14'b01111011011111:	sigmoid = 21'b111111111111111111111;
		14'b01111011100000:	sigmoid = 21'b111111111111111111111;
		14'b01111011100001:	sigmoid = 21'b111111111111111111111;
		14'b01111011100010:	sigmoid = 21'b111111111111111111111;
		14'b01111011100011:	sigmoid = 21'b111111111111111111111;
		14'b01111011100100:	sigmoid = 21'b111111111111111111111;
		14'b01111011100101:	sigmoid = 21'b111111111111111111111;
		14'b01111011100110:	sigmoid = 21'b111111111111111111111;
		14'b01111011100111:	sigmoid = 21'b111111111111111111111;
		14'b01111011101000:	sigmoid = 21'b111111111111111111111;
		14'b01111011101001:	sigmoid = 21'b111111111111111111111;
		14'b01111011101010:	sigmoid = 21'b111111111111111111111;
		14'b01111011101011:	sigmoid = 21'b111111111111111111111;
		14'b01111011101100:	sigmoid = 21'b111111111111111111111;
		14'b01111011101101:	sigmoid = 21'b111111111111111111111;
		14'b01111011101110:	sigmoid = 21'b111111111111111111111;
		14'b01111011101111:	sigmoid = 21'b111111111111111111111;
		14'b01111011110000:	sigmoid = 21'b111111111111111111111;
		14'b01111011110001:	sigmoid = 21'b111111111111111111111;
		14'b01111011110010:	sigmoid = 21'b111111111111111111111;
		14'b01111011110011:	sigmoid = 21'b111111111111111111111;
		14'b01111011110100:	sigmoid = 21'b111111111111111111111;
		14'b01111011110101:	sigmoid = 21'b111111111111111111111;
		14'b01111011110110:	sigmoid = 21'b111111111111111111111;
		14'b01111011110111:	sigmoid = 21'b111111111111111111111;
		14'b01111011111000:	sigmoid = 21'b111111111111111111111;
		14'b01111011111001:	sigmoid = 21'b111111111111111111111;
		14'b01111011111010:	sigmoid = 21'b111111111111111111111;
		14'b01111011111011:	sigmoid = 21'b111111111111111111111;
		14'b01111011111100:	sigmoid = 21'b111111111111111111111;
		14'b01111011111101:	sigmoid = 21'b111111111111111111111;
		14'b01111011111110:	sigmoid = 21'b111111111111111111111;
		14'b01111011111111:	sigmoid = 21'b111111111111111111111;
		14'b01111100000000:	sigmoid = 21'b111111111111111111111;
		14'b01111100000001:	sigmoid = 21'b111111111111111111111;
		14'b01111100000010:	sigmoid = 21'b111111111111111111111;
		14'b01111100000011:	sigmoid = 21'b111111111111111111111;
		14'b01111100000100:	sigmoid = 21'b111111111111111111111;
		14'b01111100000101:	sigmoid = 21'b111111111111111111111;
		14'b01111100000110:	sigmoid = 21'b111111111111111111111;
		14'b01111100000111:	sigmoid = 21'b111111111111111111111;
		14'b01111100001000:	sigmoid = 21'b111111111111111111111;
		14'b01111100001001:	sigmoid = 21'b111111111111111111111;
		14'b01111100001010:	sigmoid = 21'b111111111111111111111;
		14'b01111100001011:	sigmoid = 21'b111111111111111111111;
		14'b01111100001100:	sigmoid = 21'b111111111111111111111;
		14'b01111100001101:	sigmoid = 21'b111111111111111111111;
		14'b01111100001110:	sigmoid = 21'b111111111111111111111;
		14'b01111100001111:	sigmoid = 21'b111111111111111111111;
		14'b01111100010000:	sigmoid = 21'b111111111111111111111;
		14'b01111100010001:	sigmoid = 21'b111111111111111111111;
		14'b01111100010010:	sigmoid = 21'b111111111111111111111;
		14'b01111100010011:	sigmoid = 21'b111111111111111111111;
		14'b01111100010100:	sigmoid = 21'b111111111111111111111;
		14'b01111100010101:	sigmoid = 21'b111111111111111111111;
		14'b01111100010110:	sigmoid = 21'b111111111111111111111;
		14'b01111100010111:	sigmoid = 21'b111111111111111111111;
		14'b01111100011000:	sigmoid = 21'b111111111111111111111;
		14'b01111100011001:	sigmoid = 21'b111111111111111111111;
		14'b01111100011010:	sigmoid = 21'b111111111111111111111;
		14'b01111100011011:	sigmoid = 21'b111111111111111111111;
		14'b01111100011100:	sigmoid = 21'b111111111111111111111;
		14'b01111100011101:	sigmoid = 21'b111111111111111111111;
		14'b01111100011110:	sigmoid = 21'b111111111111111111111;
		14'b01111100011111:	sigmoid = 21'b111111111111111111111;
		14'b01111100100000:	sigmoid = 21'b111111111111111111111;
		14'b01111100100001:	sigmoid = 21'b111111111111111111111;
		14'b01111100100010:	sigmoid = 21'b111111111111111111111;
		14'b01111100100011:	sigmoid = 21'b111111111111111111111;
		14'b01111100100100:	sigmoid = 21'b111111111111111111111;
		14'b01111100100101:	sigmoid = 21'b111111111111111111111;
		14'b01111100100110:	sigmoid = 21'b111111111111111111111;
		14'b01111100100111:	sigmoid = 21'b111111111111111111111;
		14'b01111100101000:	sigmoid = 21'b111111111111111111111;
		14'b01111100101001:	sigmoid = 21'b111111111111111111111;
		14'b01111100101010:	sigmoid = 21'b111111111111111111111;
		14'b01111100101011:	sigmoid = 21'b111111111111111111111;
		14'b01111100101100:	sigmoid = 21'b111111111111111111111;
		14'b01111100101101:	sigmoid = 21'b111111111111111111111;
		14'b01111100101110:	sigmoid = 21'b111111111111111111111;
		14'b01111100101111:	sigmoid = 21'b111111111111111111111;
		14'b01111100110000:	sigmoid = 21'b111111111111111111111;
		14'b01111100110001:	sigmoid = 21'b111111111111111111111;
		14'b01111100110010:	sigmoid = 21'b111111111111111111111;
		14'b01111100110011:	sigmoid = 21'b111111111111111111111;
		14'b01111100110100:	sigmoid = 21'b111111111111111111111;
		14'b01111100110101:	sigmoid = 21'b111111111111111111111;
		14'b01111100110110:	sigmoid = 21'b111111111111111111111;
		14'b01111100110111:	sigmoid = 21'b111111111111111111111;
		14'b01111100111000:	sigmoid = 21'b111111111111111111111;
		14'b01111100111001:	sigmoid = 21'b111111111111111111111;
		14'b01111100111010:	sigmoid = 21'b111111111111111111111;
		14'b01111100111011:	sigmoid = 21'b111111111111111111111;
		14'b01111100111100:	sigmoid = 21'b111111111111111111111;
		14'b01111100111101:	sigmoid = 21'b111111111111111111111;
		14'b01111100111110:	sigmoid = 21'b111111111111111111111;
		14'b01111100111111:	sigmoid = 21'b111111111111111111111;
		14'b01111101000000:	sigmoid = 21'b111111111111111111111;
		14'b01111101000001:	sigmoid = 21'b111111111111111111111;
		14'b01111101000010:	sigmoid = 21'b111111111111111111111;
		14'b01111101000011:	sigmoid = 21'b111111111111111111111;
		14'b01111101000100:	sigmoid = 21'b111111111111111111111;
		14'b01111101000101:	sigmoid = 21'b111111111111111111111;
		14'b01111101000110:	sigmoid = 21'b111111111111111111111;
		14'b01111101000111:	sigmoid = 21'b111111111111111111111;
		14'b01111101001000:	sigmoid = 21'b111111111111111111111;
		14'b01111101001001:	sigmoid = 21'b111111111111111111111;
		14'b01111101001010:	sigmoid = 21'b111111111111111111111;
		14'b01111101001011:	sigmoid = 21'b111111111111111111111;
		14'b01111101001100:	sigmoid = 21'b111111111111111111111;
		14'b01111101001101:	sigmoid = 21'b111111111111111111111;
		14'b01111101001110:	sigmoid = 21'b111111111111111111111;
		14'b01111101001111:	sigmoid = 21'b111111111111111111111;
		14'b01111101010000:	sigmoid = 21'b111111111111111111111;
		14'b01111101010001:	sigmoid = 21'b111111111111111111111;
		14'b01111101010010:	sigmoid = 21'b111111111111111111111;
		14'b01111101010011:	sigmoid = 21'b111111111111111111111;
		14'b01111101010100:	sigmoid = 21'b111111111111111111111;
		14'b01111101010101:	sigmoid = 21'b111111111111111111111;
		14'b01111101010110:	sigmoid = 21'b111111111111111111111;
		14'b01111101010111:	sigmoid = 21'b111111111111111111111;
		14'b01111101011000:	sigmoid = 21'b111111111111111111111;
		14'b01111101011001:	sigmoid = 21'b111111111111111111111;
		14'b01111101011010:	sigmoid = 21'b111111111111111111111;
		14'b01111101011011:	sigmoid = 21'b111111111111111111111;
		14'b01111101011100:	sigmoid = 21'b111111111111111111111;
		14'b01111101011101:	sigmoid = 21'b111111111111111111111;
		14'b01111101011110:	sigmoid = 21'b111111111111111111111;
		14'b01111101011111:	sigmoid = 21'b111111111111111111111;
		14'b01111101100000:	sigmoid = 21'b111111111111111111111;
		14'b01111101100001:	sigmoid = 21'b111111111111111111111;
		14'b01111101100010:	sigmoid = 21'b111111111111111111111;
		14'b01111101100011:	sigmoid = 21'b111111111111111111111;
		14'b01111101100100:	sigmoid = 21'b111111111111111111111;
		14'b01111101100101:	sigmoid = 21'b111111111111111111111;
		14'b01111101100110:	sigmoid = 21'b111111111111111111111;
		14'b01111101100111:	sigmoid = 21'b111111111111111111111;
		14'b01111101101000:	sigmoid = 21'b111111111111111111111;
		14'b01111101101001:	sigmoid = 21'b111111111111111111111;
		14'b01111101101010:	sigmoid = 21'b111111111111111111111;
		14'b01111101101011:	sigmoid = 21'b111111111111111111111;
		14'b01111101101100:	sigmoid = 21'b111111111111111111111;
		14'b01111101101101:	sigmoid = 21'b111111111111111111111;
		14'b01111101101110:	sigmoid = 21'b111111111111111111111;
		14'b01111101101111:	sigmoid = 21'b111111111111111111111;
		14'b01111101110000:	sigmoid = 21'b111111111111111111111;
		14'b01111101110001:	sigmoid = 21'b111111111111111111111;
		14'b01111101110010:	sigmoid = 21'b111111111111111111111;
		14'b01111101110011:	sigmoid = 21'b111111111111111111111;
		14'b01111101110100:	sigmoid = 21'b111111111111111111111;
		14'b01111101110101:	sigmoid = 21'b111111111111111111111;
		14'b01111101110110:	sigmoid = 21'b111111111111111111111;
		14'b01111101110111:	sigmoid = 21'b111111111111111111111;
		14'b01111101111000:	sigmoid = 21'b111111111111111111111;
		14'b01111101111001:	sigmoid = 21'b111111111111111111111;
		14'b01111101111010:	sigmoid = 21'b111111111111111111111;
		14'b01111101111011:	sigmoid = 21'b111111111111111111111;
		14'b01111101111100:	sigmoid = 21'b111111111111111111111;
		14'b01111101111101:	sigmoid = 21'b111111111111111111111;
		14'b01111101111110:	sigmoid = 21'b111111111111111111111;
		14'b01111101111111:	sigmoid = 21'b111111111111111111111;
		14'b01111110000000:	sigmoid = 21'b111111111111111111111;
		14'b01111110000001:	sigmoid = 21'b111111111111111111111;
		14'b01111110000010:	sigmoid = 21'b111111111111111111111;
		14'b01111110000011:	sigmoid = 21'b111111111111111111111;
		14'b01111110000100:	sigmoid = 21'b111111111111111111111;
		14'b01111110000101:	sigmoid = 21'b111111111111111111111;
		14'b01111110000110:	sigmoid = 21'b111111111111111111111;
		14'b01111110000111:	sigmoid = 21'b111111111111111111111;
		14'b01111110001000:	sigmoid = 21'b111111111111111111111;
		14'b01111110001001:	sigmoid = 21'b111111111111111111111;
		14'b01111110001010:	sigmoid = 21'b111111111111111111111;
		14'b01111110001011:	sigmoid = 21'b111111111111111111111;
		14'b01111110001100:	sigmoid = 21'b111111111111111111111;
		14'b01111110001101:	sigmoid = 21'b111111111111111111111;
		14'b01111110001110:	sigmoid = 21'b111111111111111111111;
		14'b01111110001111:	sigmoid = 21'b111111111111111111111;
		14'b01111110010000:	sigmoid = 21'b111111111111111111111;
		14'b01111110010001:	sigmoid = 21'b111111111111111111111;
		14'b01111110010010:	sigmoid = 21'b111111111111111111111;
		14'b01111110010011:	sigmoid = 21'b111111111111111111111;
		14'b01111110010100:	sigmoid = 21'b111111111111111111111;
		14'b01111110010101:	sigmoid = 21'b111111111111111111111;
		14'b01111110010110:	sigmoid = 21'b111111111111111111111;
		14'b01111110010111:	sigmoid = 21'b111111111111111111111;
		14'b01111110011000:	sigmoid = 21'b111111111111111111111;
		14'b01111110011001:	sigmoid = 21'b111111111111111111111;
		14'b01111110011010:	sigmoid = 21'b111111111111111111111;
		14'b01111110011011:	sigmoid = 21'b111111111111111111111;
		14'b01111110011100:	sigmoid = 21'b111111111111111111111;
		14'b01111110011101:	sigmoid = 21'b111111111111111111111;
		14'b01111110011110:	sigmoid = 21'b111111111111111111111;
		14'b01111110011111:	sigmoid = 21'b111111111111111111111;
		14'b01111110100000:	sigmoid = 21'b111111111111111111111;
		14'b01111110100001:	sigmoid = 21'b111111111111111111111;
		14'b01111110100010:	sigmoid = 21'b111111111111111111111;
		14'b01111110100011:	sigmoid = 21'b111111111111111111111;
		14'b01111110100100:	sigmoid = 21'b111111111111111111111;
		14'b01111110100101:	sigmoid = 21'b111111111111111111111;
		14'b01111110100110:	sigmoid = 21'b111111111111111111111;
		14'b01111110100111:	sigmoid = 21'b111111111111111111111;
		14'b01111110101000:	sigmoid = 21'b111111111111111111111;
		14'b01111110101001:	sigmoid = 21'b111111111111111111111;
		14'b01111110101010:	sigmoid = 21'b111111111111111111111;
		14'b01111110101011:	sigmoid = 21'b111111111111111111111;
		14'b01111110101100:	sigmoid = 21'b111111111111111111111;
		14'b01111110101101:	sigmoid = 21'b111111111111111111111;
		14'b01111110101110:	sigmoid = 21'b111111111111111111111;
		14'b01111110101111:	sigmoid = 21'b111111111111111111111;
		14'b01111110110000:	sigmoid = 21'b111111111111111111111;
		14'b01111110110001:	sigmoid = 21'b111111111111111111111;
		14'b01111110110010:	sigmoid = 21'b111111111111111111111;
		14'b01111110110011:	sigmoid = 21'b111111111111111111111;
		14'b01111110110100:	sigmoid = 21'b111111111111111111111;
		14'b01111110110101:	sigmoid = 21'b111111111111111111111;
		14'b01111110110110:	sigmoid = 21'b111111111111111111111;
		14'b01111110110111:	sigmoid = 21'b111111111111111111111;
		14'b01111110111000:	sigmoid = 21'b111111111111111111111;
		14'b01111110111001:	sigmoid = 21'b111111111111111111111;
		14'b01111110111010:	sigmoid = 21'b111111111111111111111;
		14'b01111110111011:	sigmoid = 21'b111111111111111111111;
		14'b01111110111100:	sigmoid = 21'b111111111111111111111;
		14'b01111110111101:	sigmoid = 21'b111111111111111111111;
		14'b01111110111110:	sigmoid = 21'b111111111111111111111;
		14'b01111110111111:	sigmoid = 21'b111111111111111111111;
		14'b01111111000000:	sigmoid = 21'b111111111111111111111;
		14'b01111111000001:	sigmoid = 21'b111111111111111111111;
		14'b01111111000010:	sigmoid = 21'b111111111111111111111;
		14'b01111111000011:	sigmoid = 21'b111111111111111111111;
		14'b01111111000100:	sigmoid = 21'b111111111111111111111;
		14'b01111111000101:	sigmoid = 21'b111111111111111111111;
		14'b01111111000110:	sigmoid = 21'b111111111111111111111;
		14'b01111111000111:	sigmoid = 21'b111111111111111111111;
		14'b01111111001000:	sigmoid = 21'b111111111111111111111;
		14'b01111111001001:	sigmoid = 21'b111111111111111111111;
		14'b01111111001010:	sigmoid = 21'b111111111111111111111;
		14'b01111111001011:	sigmoid = 21'b111111111111111111111;
		14'b01111111001100:	sigmoid = 21'b111111111111111111111;
		14'b01111111001101:	sigmoid = 21'b111111111111111111111;
		14'b01111111001110:	sigmoid = 21'b111111111111111111111;
		14'b01111111001111:	sigmoid = 21'b111111111111111111111;
		14'b01111111010000:	sigmoid = 21'b111111111111111111111;
		14'b01111111010001:	sigmoid = 21'b111111111111111111111;
		14'b01111111010010:	sigmoid = 21'b111111111111111111111;
		14'b01111111010011:	sigmoid = 21'b111111111111111111111;
		14'b01111111010100:	sigmoid = 21'b111111111111111111111;
		14'b01111111010101:	sigmoid = 21'b111111111111111111111;
		14'b01111111010110:	sigmoid = 21'b111111111111111111111;
		14'b01111111010111:	sigmoid = 21'b111111111111111111111;
		14'b01111111011000:	sigmoid = 21'b111111111111111111111;
		14'b01111111011001:	sigmoid = 21'b111111111111111111111;
		14'b01111111011010:	sigmoid = 21'b111111111111111111111;
		14'b01111111011011:	sigmoid = 21'b111111111111111111111;
		14'b01111111011100:	sigmoid = 21'b111111111111111111111;
		14'b01111111011101:	sigmoid = 21'b111111111111111111111;
		14'b01111111011110:	sigmoid = 21'b111111111111111111111;
		14'b01111111011111:	sigmoid = 21'b111111111111111111111;
		14'b01111111100000:	sigmoid = 21'b111111111111111111111;
		14'b01111111100001:	sigmoid = 21'b111111111111111111111;
		14'b01111111100010:	sigmoid = 21'b111111111111111111111;
		14'b01111111100011:	sigmoid = 21'b111111111111111111111;
		14'b01111111100100:	sigmoid = 21'b111111111111111111111;
		14'b01111111100101:	sigmoid = 21'b111111111111111111111;
		14'b01111111100110:	sigmoid = 21'b111111111111111111111;
		14'b01111111100111:	sigmoid = 21'b111111111111111111111;
		14'b01111111101000:	sigmoid = 21'b111111111111111111111;
		14'b01111111101001:	sigmoid = 21'b111111111111111111111;
		14'b01111111101010:	sigmoid = 21'b111111111111111111111;
		14'b01111111101011:	sigmoid = 21'b111111111111111111111;
		14'b01111111101100:	sigmoid = 21'b111111111111111111111;
		14'b01111111101101:	sigmoid = 21'b111111111111111111111;
		14'b01111111101110:	sigmoid = 21'b111111111111111111111;
		14'b01111111101111:	sigmoid = 21'b111111111111111111111;
		14'b01111111110000:	sigmoid = 21'b111111111111111111111;
		14'b01111111110001:	sigmoid = 21'b111111111111111111111;
		14'b01111111110010:	sigmoid = 21'b111111111111111111111;
		14'b01111111110011:	sigmoid = 21'b111111111111111111111;
		14'b01111111110100:	sigmoid = 21'b111111111111111111111;
		14'b01111111110101:	sigmoid = 21'b111111111111111111111;
		14'b01111111110110:	sigmoid = 21'b111111111111111111111;
		14'b01111111110111:	sigmoid = 21'b111111111111111111111;
		14'b01111111111000:	sigmoid = 21'b111111111111111111111;
		14'b01111111111001:	sigmoid = 21'b111111111111111111111;
		14'b01111111111010:	sigmoid = 21'b111111111111111111111;
		14'b01111111111011:	sigmoid = 21'b111111111111111111111;
		14'b01111111111100:	sigmoid = 21'b111111111111111111111;
		14'b01111111111101:	sigmoid = 21'b111111111111111111111;
		14'b01111111111110:	sigmoid = 21'b111111111111111111111;
		14'b01111111111111:	sigmoid = 21'b111111111111111111111;

	endcase
endmodule

// __________________________________________________________________________________________________________ //
// __________________________________________________________________________________________________________ //

/*  SIGMOID PRIME TABLE:
	Original z = 16b = 1,5,10 => -32 to +32
	Domain z used here = 10b = 1,3,6 => -8 to +8, 0.015625 precision. These are bits [13:4] of original z
	When z<-8 or z>8, f'(z)=0. When z=0, f'(z)=0.25
	Range f'(z) = 8b = 0,-2,10 => 0 to 0.25, 0.0009766 precision.
	Final sigmoid output value = 16b = 1,5,10. DIFFERENT FROM SIGMOID: 8 MSB are all 0. Bits [7:0] of final value are calculated f'(z) */
module sig_prime #(
	parameter width = 32, 
	parameter int_bits = 10,
	parameter frac_bits = 21
)(
	input clk,
	input [width-1:0] z,
	output reg[width-1:0] sp_out
);
	
	reg [17:0] sigmoid_prime;
	/*real real_z, real_sp;

	

	always @(posedge clk)begin
		real_z = z/2**(frac_bits)-z[width-1]*2.0**(1+int_bits);
		real_sp = 1.0/(1+2.71828**(-real_z))*(1.0-1.0/(1+2.71828**(-real_z)));
		sp_out = real_sp*2**(frac_bits)+10;
	end*/
	always @(posedge clk)
	sp_out = (z[width-1:width-int_bits+2] == 0 ||&z[width-1:width-int_bits+2])? 
			{{(int_bits+2){1'b0}},sigmoid_prime}:1;
	// If condition is not met, z is too high or too low. In that case, f'(z)=0

	always @(z[frac_bits+4:frac_bits-9])
	case (z[frac_bits+4:frac_bits-9])
		//sign, 3bits_i, 6bits_f ~ 0.015625  --->   8bits_f ~ 0.0009766(3~10)
		14'b10000000000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000000111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000001111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000010111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000011111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000100111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000101111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000110111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10000111111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001000111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001001111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001010111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001011111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001100111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001101111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001110111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10001111111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010000111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010001111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010010111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010011111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010100111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010101111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010110111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10010111111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011000111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011001111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011010111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011011111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011100111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011101111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011110111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10011111111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000101111:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000110000:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000110001:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000110010:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000110011:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000110100:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000110101:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000110110:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000110111:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000111000:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000111001:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000111010:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000111011:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000111100:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000111101:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000111110:	sigmoid_prime = 18'b000000000000000001;
		14'b10100000111111:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001000000:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001000001:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001000010:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001000011:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001000100:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001000101:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001000110:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001000111:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001001000:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001001001:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001001010:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001001011:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001001100:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001001101:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001001110:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001001111:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001010000:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001010001:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001010010:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001010011:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001010100:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001010101:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001010110:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001010111:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001011000:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001011001:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001011010:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001011011:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001011100:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001011101:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001011110:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001011111:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001100000:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001100001:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001100010:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001100011:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001100100:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001100101:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001100110:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001100111:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001101000:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001101001:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001101010:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001101011:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001101100:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001101101:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001101110:	sigmoid_prime = 18'b000000000000000001;
		14'b10100001101111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001110000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001110001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001110010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001110011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001110100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001110101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001110110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001110111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001111000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001111001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001111010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001111011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001111100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001111101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001111110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100001111111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010000000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010000001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010000010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010000011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010000100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010000101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010000110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010000111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010001000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010001001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010001010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010001011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010001100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010001101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010001110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010001111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010010000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010010001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010010010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010010011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010010100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010010101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010010110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010010111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010011000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010011001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010011010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010011011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010011100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010011101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010011110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010011111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010100000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010100001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010100010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010100011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010100100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010100101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010100110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010100111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010101000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010101001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010101010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010101011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010101100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010101101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010101110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010101111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010110000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010110001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010110010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010110011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010110100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010110101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010110110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010110111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010111000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010111001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010111010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010111011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010111100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010111101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010111110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100010111111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011000000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011000001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011000010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011000011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011000100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011000101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011000110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011000111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011001000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011001001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011001010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011001011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011001100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011001101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011001110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011001111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011010000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011010001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011010010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011010011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011010100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011010101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011010110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011010111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011011000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011011001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011011010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011011011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011011100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011011101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011011110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011011111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011100000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011100001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011100010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011100011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011100100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011100101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011100110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011100111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011101000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011101001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011101010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011101011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011101100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011101101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011101110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011101111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011110000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011110001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011110010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011110011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011110100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011110101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011110110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011110111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011111000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011111001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011111010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011111011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011111100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011111101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011111110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100011111111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100000000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100000001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100000010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100000011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100000100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100000101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100000110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100000111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100001000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100001001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100001010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100001011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100001100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100001101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100001110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100001111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100010000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100010001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100010010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100010011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100010100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100010101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100010110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100010111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100011000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100011001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100011010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100011011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100011100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100011101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100011110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100011111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100100000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100100001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100100010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100100011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100100100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100100101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100100110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100100111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100101000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100101001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100101010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100101011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100101100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100101101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100101110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100101111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100110000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100110001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100110010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100110011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100110100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100110101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100110110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100110111:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100111000:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100111001:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100111010:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100111011:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100111100:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100111101:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100111110:	sigmoid_prime = 18'b000000000000000010;
		14'b10100100111111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101000000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101000001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101000010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101000011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101000100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101000101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101000110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101000111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101001000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101001001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101001010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101001011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101001100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101001101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101001110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101001111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101010000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101010001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101010010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101010011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101010100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101010101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101010110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101010111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101011000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101011001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101011010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101011011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101011100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101011101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101011110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101011111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101100000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101100001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101100010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101100011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101100100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101100101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101100110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101100111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101101000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101101001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101101010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101101011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101101100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101101101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101101110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101101111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101110000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101110001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101110010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101110011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101110100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101110101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101110110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101110111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101111000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101111001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101111010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101111011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101111100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101111101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101111110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100101111111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110000000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110000001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110000010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110000011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110000100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110000101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110000110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110000111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110001000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110001001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110001010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110001011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110001100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110001101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110001110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110001111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110010000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110010001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110010010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110010011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110010100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110010101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110010110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110010111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110011000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110011001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110011010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110011011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110011100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110011101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110011110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110011111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110100000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110100001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110100010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110100011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110100100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110100101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110100110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110100111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110101000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110101001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110101010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110101011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110101100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110101101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110101110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110101111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110110000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110110001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110110010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110110011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110110100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110110101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110110110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110110111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110111000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110111001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110111010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110111011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110111100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110111101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110111110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100110111111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111000000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111000001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111000010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111000011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111000100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111000101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111000110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111000111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111001000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111001001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111001010:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111001011:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111001100:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111001101:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111001110:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111001111:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111010000:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111010001:	sigmoid_prime = 18'b000000000000000011;
		14'b10100111010010:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111010011:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111010100:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111010101:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111010110:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111010111:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111011000:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111011001:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111011010:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111011011:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111011100:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111011101:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111011110:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111011111:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111100000:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111100001:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111100010:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111100011:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111100100:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111100101:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111100110:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111100111:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111101000:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111101001:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111101010:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111101011:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111101100:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111101101:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111101110:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111101111:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111110000:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111110001:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111110010:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111110011:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111110100:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111110101:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111110110:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111110111:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111111000:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111111001:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111111010:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111111011:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111111100:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111111101:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111111110:	sigmoid_prime = 18'b000000000000000100;
		14'b10100111111111:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000000000:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000000001:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000000010:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000000011:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000000100:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000000101:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000000110:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000000111:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000001000:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000001001:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000001010:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000001011:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000001100:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000001101:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000001110:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000001111:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000010000:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000010001:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000010010:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000010011:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000010100:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000010101:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000010110:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000010111:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000011000:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000011001:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000011010:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000011011:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000011100:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000011101:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000011110:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000011111:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000100000:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000100001:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000100010:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000100011:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000100100:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000100101:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000100110:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000100111:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000101000:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000101001:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000101010:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000101011:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000101100:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000101101:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000101110:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000101111:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000110000:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000110001:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000110010:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000110011:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000110100:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000110101:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000110110:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000110111:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000111000:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000111001:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000111010:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000111011:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000111100:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000111101:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000111110:	sigmoid_prime = 18'b000000000000000100;
		14'b10101000111111:	sigmoid_prime = 18'b000000000000000100;
		14'b10101001000000:	sigmoid_prime = 18'b000000000000000100;
		14'b10101001000001:	sigmoid_prime = 18'b000000000000000100;
		14'b10101001000010:	sigmoid_prime = 18'b000000000000000100;
		14'b10101001000011:	sigmoid_prime = 18'b000000000000000100;
		14'b10101001000100:	sigmoid_prime = 18'b000000000000000100;
		14'b10101001000101:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001000110:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001000111:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001001000:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001001001:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001001010:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001001011:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001001100:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001001101:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001001110:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001001111:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001010000:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001010001:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001010010:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001010011:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001010100:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001010101:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001010110:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001010111:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001011000:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001011001:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001011010:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001011011:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001011100:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001011101:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001011110:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001011111:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001100000:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001100001:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001100010:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001100011:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001100100:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001100101:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001100110:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001100111:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001101000:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001101001:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001101010:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001101011:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001101100:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001101101:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001101110:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001101111:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001110000:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001110001:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001110010:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001110011:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001110100:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001110101:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001110110:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001110111:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001111000:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001111001:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001111010:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001111011:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001111100:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001111101:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001111110:	sigmoid_prime = 18'b000000000000000101;
		14'b10101001111111:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010000000:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010000001:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010000010:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010000011:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010000100:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010000101:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010000110:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010000111:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010001000:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010001001:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010001010:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010001011:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010001100:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010001101:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010001110:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010001111:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010010000:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010010001:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010010010:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010010011:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010010100:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010010101:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010010110:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010010111:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010011000:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010011001:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010011010:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010011011:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010011100:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010011101:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010011110:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010011111:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010100000:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010100001:	sigmoid_prime = 18'b000000000000000101;
		14'b10101010100010:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010100011:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010100100:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010100101:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010100110:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010100111:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010101000:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010101001:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010101010:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010101011:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010101100:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010101101:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010101110:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010101111:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010110000:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010110001:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010110010:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010110011:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010110100:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010110101:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010110110:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010110111:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010111000:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010111001:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010111010:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010111011:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010111100:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010111101:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010111110:	sigmoid_prime = 18'b000000000000000110;
		14'b10101010111111:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011000000:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011000001:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011000010:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011000011:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011000100:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011000101:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011000110:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011000111:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011001000:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011001001:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011001010:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011001011:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011001100:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011001101:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011001110:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011001111:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011010000:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011010001:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011010010:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011010011:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011010100:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011010101:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011010110:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011010111:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011011000:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011011001:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011011010:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011011011:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011011100:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011011101:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011011110:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011011111:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011100000:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011100001:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011100010:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011100011:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011100100:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011100101:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011100110:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011100111:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011101000:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011101001:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011101010:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011101011:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011101100:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011101101:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011101110:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011101111:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011110000:	sigmoid_prime = 18'b000000000000000110;
		14'b10101011110001:	sigmoid_prime = 18'b000000000000000111;
		14'b10101011110010:	sigmoid_prime = 18'b000000000000000111;
		14'b10101011110011:	sigmoid_prime = 18'b000000000000000111;
		14'b10101011110100:	sigmoid_prime = 18'b000000000000000111;
		14'b10101011110101:	sigmoid_prime = 18'b000000000000000111;
		14'b10101011110110:	sigmoid_prime = 18'b000000000000000111;
		14'b10101011110111:	sigmoid_prime = 18'b000000000000000111;
		14'b10101011111000:	sigmoid_prime = 18'b000000000000000111;
		14'b10101011111001:	sigmoid_prime = 18'b000000000000000111;
		14'b10101011111010:	sigmoid_prime = 18'b000000000000000111;
		14'b10101011111011:	sigmoid_prime = 18'b000000000000000111;
		14'b10101011111100:	sigmoid_prime = 18'b000000000000000111;
		14'b10101011111101:	sigmoid_prime = 18'b000000000000000111;
		14'b10101011111110:	sigmoid_prime = 18'b000000000000000111;
		14'b10101011111111:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100000000:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100000001:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100000010:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100000011:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100000100:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100000101:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100000110:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100000111:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100001000:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100001001:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100001010:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100001011:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100001100:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100001101:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100001110:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100001111:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100010000:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100010001:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100010010:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100010011:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100010100:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100010101:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100010110:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100010111:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100011000:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100011001:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100011010:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100011011:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100011100:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100011101:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100011110:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100011111:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100100000:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100100001:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100100010:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100100011:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100100100:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100100101:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100100110:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100100111:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100101000:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100101001:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100101010:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100101011:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100101100:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100101101:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100101110:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100101111:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100110000:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100110001:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100110010:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100110011:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100110100:	sigmoid_prime = 18'b000000000000000111;
		14'b10101100110101:	sigmoid_prime = 18'b000000000000001000;
		14'b10101100110110:	sigmoid_prime = 18'b000000000000001000;
		14'b10101100110111:	sigmoid_prime = 18'b000000000000001000;
		14'b10101100111000:	sigmoid_prime = 18'b000000000000001000;
		14'b10101100111001:	sigmoid_prime = 18'b000000000000001000;
		14'b10101100111010:	sigmoid_prime = 18'b000000000000001000;
		14'b10101100111011:	sigmoid_prime = 18'b000000000000001000;
		14'b10101100111100:	sigmoid_prime = 18'b000000000000001000;
		14'b10101100111101:	sigmoid_prime = 18'b000000000000001000;
		14'b10101100111110:	sigmoid_prime = 18'b000000000000001000;
		14'b10101100111111:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101000000:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101000001:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101000010:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101000011:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101000100:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101000101:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101000110:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101000111:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101001000:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101001001:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101001010:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101001011:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101001100:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101001101:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101001110:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101001111:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101010000:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101010001:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101010010:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101010011:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101010100:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101010101:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101010110:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101010111:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101011000:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101011001:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101011010:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101011011:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101011100:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101011101:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101011110:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101011111:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101100000:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101100001:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101100010:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101100011:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101100100:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101100101:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101100110:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101100111:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101101000:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101101001:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101101010:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101101011:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101101100:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101101101:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101101110:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101101111:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101110000:	sigmoid_prime = 18'b000000000000001000;
		14'b10101101110001:	sigmoid_prime = 18'b000000000000001001;
		14'b10101101110010:	sigmoid_prime = 18'b000000000000001001;
		14'b10101101110011:	sigmoid_prime = 18'b000000000000001001;
		14'b10101101110100:	sigmoid_prime = 18'b000000000000001001;
		14'b10101101110101:	sigmoid_prime = 18'b000000000000001001;
		14'b10101101110110:	sigmoid_prime = 18'b000000000000001001;
		14'b10101101110111:	sigmoid_prime = 18'b000000000000001001;
		14'b10101101111000:	sigmoid_prime = 18'b000000000000001001;
		14'b10101101111001:	sigmoid_prime = 18'b000000000000001001;
		14'b10101101111010:	sigmoid_prime = 18'b000000000000001001;
		14'b10101101111011:	sigmoid_prime = 18'b000000000000001001;
		14'b10101101111100:	sigmoid_prime = 18'b000000000000001001;
		14'b10101101111101:	sigmoid_prime = 18'b000000000000001001;
		14'b10101101111110:	sigmoid_prime = 18'b000000000000001001;
		14'b10101101111111:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110000000:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110000001:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110000010:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110000011:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110000100:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110000101:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110000110:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110000111:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110001000:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110001001:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110001010:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110001011:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110001100:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110001101:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110001110:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110001111:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110010000:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110010001:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110010010:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110010011:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110010100:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110010101:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110010110:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110010111:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110011000:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110011001:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110011010:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110011011:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110011100:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110011101:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110011110:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110011111:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110100000:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110100001:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110100010:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110100011:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110100100:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110100101:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110100110:	sigmoid_prime = 18'b000000000000001001;
		14'b10101110100111:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110101000:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110101001:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110101010:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110101011:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110101100:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110101101:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110101110:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110101111:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110110000:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110110001:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110110010:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110110011:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110110100:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110110101:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110110110:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110110111:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110111000:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110111001:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110111010:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110111011:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110111100:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110111101:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110111110:	sigmoid_prime = 18'b000000000000001010;
		14'b10101110111111:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111000000:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111000001:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111000010:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111000011:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111000100:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111000101:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111000110:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111000111:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111001000:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111001001:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111001010:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111001011:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111001100:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111001101:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111001110:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111001111:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111010000:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111010001:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111010010:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111010011:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111010100:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111010101:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111010110:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111010111:	sigmoid_prime = 18'b000000000000001010;
		14'b10101111011000:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111011001:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111011010:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111011011:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111011100:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111011101:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111011110:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111011111:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111100000:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111100001:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111100010:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111100011:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111100100:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111100101:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111100110:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111100111:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111101000:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111101001:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111101010:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111101011:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111101100:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111101101:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111101110:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111101111:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111110000:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111110001:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111110010:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111110011:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111110100:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111110101:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111110110:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111110111:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111111000:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111111001:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111111010:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111111011:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111111100:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111111101:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111111110:	sigmoid_prime = 18'b000000000000001011;
		14'b10101111111111:	sigmoid_prime = 18'b000000000000001011;
		14'b10110000000000:	sigmoid_prime = 18'b000000000000001011;
		14'b10110000000001:	sigmoid_prime = 18'b000000000000001011;
		14'b10110000000010:	sigmoid_prime = 18'b000000000000001011;
		14'b10110000000011:	sigmoid_prime = 18'b000000000000001011;
		14'b10110000000100:	sigmoid_prime = 18'b000000000000001011;
		14'b10110000000101:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000000110:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000000111:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000001000:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000001001:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000001010:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000001011:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000001100:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000001101:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000001110:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000001111:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000010000:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000010001:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000010010:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000010011:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000010100:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000010101:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000010110:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000010111:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000011000:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000011001:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000011010:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000011011:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000011100:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000011101:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000011110:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000011111:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000100000:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000100001:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000100010:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000100011:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000100100:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000100101:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000100110:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000100111:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000101000:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000101001:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000101010:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000101011:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000101100:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000101101:	sigmoid_prime = 18'b000000000000001100;
		14'b10110000101110:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000101111:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000110000:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000110001:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000110010:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000110011:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000110100:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000110101:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000110110:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000110111:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000111000:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000111001:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000111010:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000111011:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000111100:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000111101:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000111110:	sigmoid_prime = 18'b000000000000001101;
		14'b10110000111111:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001000000:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001000001:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001000010:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001000011:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001000100:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001000101:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001000110:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001000111:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001001000:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001001001:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001001010:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001001011:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001001100:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001001101:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001001110:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001001111:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001010000:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001010001:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001010010:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001010011:	sigmoid_prime = 18'b000000000000001101;
		14'b10110001010100:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001010101:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001010110:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001010111:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001011000:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001011001:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001011010:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001011011:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001011100:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001011101:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001011110:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001011111:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001100000:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001100001:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001100010:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001100011:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001100100:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001100101:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001100110:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001100111:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001101000:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001101001:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001101010:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001101011:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001101100:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001101101:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001101110:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001101111:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001110000:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001110001:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001110010:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001110011:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001110100:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001110101:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001110110:	sigmoid_prime = 18'b000000000000001110;
		14'b10110001110111:	sigmoid_prime = 18'b000000000000001111;
		14'b10110001111000:	sigmoid_prime = 18'b000000000000001111;
		14'b10110001111001:	sigmoid_prime = 18'b000000000000001111;
		14'b10110001111010:	sigmoid_prime = 18'b000000000000001111;
		14'b10110001111011:	sigmoid_prime = 18'b000000000000001111;
		14'b10110001111100:	sigmoid_prime = 18'b000000000000001111;
		14'b10110001111101:	sigmoid_prime = 18'b000000000000001111;
		14'b10110001111110:	sigmoid_prime = 18'b000000000000001111;
		14'b10110001111111:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010000000:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010000001:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010000010:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010000011:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010000100:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010000101:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010000110:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010000111:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010001000:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010001001:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010001010:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010001011:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010001100:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010001101:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010001110:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010001111:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010010000:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010010001:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010010010:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010010011:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010010100:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010010101:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010010110:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010010111:	sigmoid_prime = 18'b000000000000001111;
		14'b10110010011000:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010011001:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010011010:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010011011:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010011100:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010011101:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010011110:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010011111:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010100000:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010100001:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010100010:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010100011:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010100100:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010100101:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010100110:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010100111:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010101000:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010101001:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010101010:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010101011:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010101100:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010101101:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010101110:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010101111:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010110000:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010110001:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010110010:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010110011:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010110100:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010110101:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010110110:	sigmoid_prime = 18'b000000000000010000;
		14'b10110010110111:	sigmoid_prime = 18'b000000000000010001;
		14'b10110010111000:	sigmoid_prime = 18'b000000000000010001;
		14'b10110010111001:	sigmoid_prime = 18'b000000000000010001;
		14'b10110010111010:	sigmoid_prime = 18'b000000000000010001;
		14'b10110010111011:	sigmoid_prime = 18'b000000000000010001;
		14'b10110010111100:	sigmoid_prime = 18'b000000000000010001;
		14'b10110010111101:	sigmoid_prime = 18'b000000000000010001;
		14'b10110010111110:	sigmoid_prime = 18'b000000000000010001;
		14'b10110010111111:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011000000:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011000001:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011000010:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011000011:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011000100:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011000101:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011000110:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011000111:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011001000:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011001001:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011001010:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011001011:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011001100:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011001101:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011001110:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011001111:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011010000:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011010001:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011010010:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011010011:	sigmoid_prime = 18'b000000000000010001;
		14'b10110011010100:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011010101:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011010110:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011010111:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011011000:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011011001:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011011010:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011011011:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011011100:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011011101:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011011110:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011011111:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011100000:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011100001:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011100010:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011100011:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011100100:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011100101:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011100110:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011100111:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011101000:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011101001:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011101010:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011101011:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011101100:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011101101:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011101110:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011101111:	sigmoid_prime = 18'b000000000000010010;
		14'b10110011110000:	sigmoid_prime = 18'b000000000000010011;
		14'b10110011110001:	sigmoid_prime = 18'b000000000000010011;
		14'b10110011110010:	sigmoid_prime = 18'b000000000000010011;
		14'b10110011110011:	sigmoid_prime = 18'b000000000000010011;
		14'b10110011110100:	sigmoid_prime = 18'b000000000000010011;
		14'b10110011110101:	sigmoid_prime = 18'b000000000000010011;
		14'b10110011110110:	sigmoid_prime = 18'b000000000000010011;
		14'b10110011110111:	sigmoid_prime = 18'b000000000000010011;
		14'b10110011111000:	sigmoid_prime = 18'b000000000000010011;
		14'b10110011111001:	sigmoid_prime = 18'b000000000000010011;
		14'b10110011111010:	sigmoid_prime = 18'b000000000000010011;
		14'b10110011111011:	sigmoid_prime = 18'b000000000000010011;
		14'b10110011111100:	sigmoid_prime = 18'b000000000000010011;
		14'b10110011111101:	sigmoid_prime = 18'b000000000000010011;
		14'b10110011111110:	sigmoid_prime = 18'b000000000000010011;
		14'b10110011111111:	sigmoid_prime = 18'b000000000000010011;
		14'b10110100000000:	sigmoid_prime = 18'b000000000000010011;
		14'b10110100000001:	sigmoid_prime = 18'b000000000000010011;
		14'b10110100000010:	sigmoid_prime = 18'b000000000000010011;
		14'b10110100000011:	sigmoid_prime = 18'b000000000000010011;
		14'b10110100000100:	sigmoid_prime = 18'b000000000000010011;
		14'b10110100000101:	sigmoid_prime = 18'b000000000000010011;
		14'b10110100000110:	sigmoid_prime = 18'b000000000000010011;
		14'b10110100000111:	sigmoid_prime = 18'b000000000000010011;
		14'b10110100001000:	sigmoid_prime = 18'b000000000000010011;
		14'b10110100001001:	sigmoid_prime = 18'b000000000000010011;
		14'b10110100001010:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100001011:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100001100:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100001101:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100001110:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100001111:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100010000:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100010001:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100010010:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100010011:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100010100:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100010101:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100010110:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100010111:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100011000:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100011001:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100011010:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100011011:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100011100:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100011101:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100011110:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100011111:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100100000:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100100001:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100100010:	sigmoid_prime = 18'b000000000000010100;
		14'b10110100100011:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100100100:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100100101:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100100110:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100100111:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100101000:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100101001:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100101010:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100101011:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100101100:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100101101:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100101110:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100101111:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100110000:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100110001:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100110010:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100110011:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100110100:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100110101:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100110110:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100110111:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100111000:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100111001:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100111010:	sigmoid_prime = 18'b000000000000010101;
		14'b10110100111011:	sigmoid_prime = 18'b000000000000010110;
		14'b10110100111100:	sigmoid_prime = 18'b000000000000010110;
		14'b10110100111101:	sigmoid_prime = 18'b000000000000010110;
		14'b10110100111110:	sigmoid_prime = 18'b000000000000010110;
		14'b10110100111111:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101000000:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101000001:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101000010:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101000011:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101000100:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101000101:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101000110:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101000111:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101001000:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101001001:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101001010:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101001011:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101001100:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101001101:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101001110:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101001111:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101010000:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101010001:	sigmoid_prime = 18'b000000000000010110;
		14'b10110101010010:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101010011:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101010100:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101010101:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101010110:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101010111:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101011000:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101011001:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101011010:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101011011:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101011100:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101011101:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101011110:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101011111:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101100000:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101100001:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101100010:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101100011:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101100100:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101100101:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101100110:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101100111:	sigmoid_prime = 18'b000000000000010111;
		14'b10110101101000:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101101001:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101101010:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101101011:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101101100:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101101101:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101101110:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101101111:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101110000:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101110001:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101110010:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101110011:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101110100:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101110101:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101110110:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101110111:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101111000:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101111001:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101111010:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101111011:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101111100:	sigmoid_prime = 18'b000000000000011000;
		14'b10110101111101:	sigmoid_prime = 18'b000000000000011001;
		14'b10110101111110:	sigmoid_prime = 18'b000000000000011001;
		14'b10110101111111:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110000000:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110000001:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110000010:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110000011:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110000100:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110000101:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110000110:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110000111:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110001000:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110001001:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110001010:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110001011:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110001100:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110001101:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110001110:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110001111:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110010000:	sigmoid_prime = 18'b000000000000011001;
		14'b10110110010001:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110010010:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110010011:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110010100:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110010101:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110010110:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110010111:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110011000:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110011001:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110011010:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110011011:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110011100:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110011101:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110011110:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110011111:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110100000:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110100001:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110100010:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110100011:	sigmoid_prime = 18'b000000000000011010;
		14'b10110110100100:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110100101:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110100110:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110100111:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110101000:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110101001:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110101010:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110101011:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110101100:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110101101:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110101110:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110101111:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110110000:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110110001:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110110010:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110110011:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110110100:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110110101:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110110110:	sigmoid_prime = 18'b000000000000011011;
		14'b10110110110111:	sigmoid_prime = 18'b000000000000011100;
		14'b10110110111000:	sigmoid_prime = 18'b000000000000011100;
		14'b10110110111001:	sigmoid_prime = 18'b000000000000011100;
		14'b10110110111010:	sigmoid_prime = 18'b000000000000011100;
		14'b10110110111011:	sigmoid_prime = 18'b000000000000011100;
		14'b10110110111100:	sigmoid_prime = 18'b000000000000011100;
		14'b10110110111101:	sigmoid_prime = 18'b000000000000011100;
		14'b10110110111110:	sigmoid_prime = 18'b000000000000011100;
		14'b10110110111111:	sigmoid_prime = 18'b000000000000011100;
		14'b10110111000000:	sigmoid_prime = 18'b000000000000011100;
		14'b10110111000001:	sigmoid_prime = 18'b000000000000011100;
		14'b10110111000010:	sigmoid_prime = 18'b000000000000011100;
		14'b10110111000011:	sigmoid_prime = 18'b000000000000011100;
		14'b10110111000100:	sigmoid_prime = 18'b000000000000011100;
		14'b10110111000101:	sigmoid_prime = 18'b000000000000011100;
		14'b10110111000110:	sigmoid_prime = 18'b000000000000011100;
		14'b10110111000111:	sigmoid_prime = 18'b000000000000011100;
		14'b10110111001000:	sigmoid_prime = 18'b000000000000011100;
		14'b10110111001001:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111001010:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111001011:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111001100:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111001101:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111001110:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111001111:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111010000:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111010001:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111010010:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111010011:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111010100:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111010101:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111010110:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111010111:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111011000:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111011001:	sigmoid_prime = 18'b000000000000011101;
		14'b10110111011010:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111011011:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111011100:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111011101:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111011110:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111011111:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111100000:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111100001:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111100010:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111100011:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111100100:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111100101:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111100110:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111100111:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111101000:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111101001:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111101010:	sigmoid_prime = 18'b000000000000011110;
		14'b10110111101011:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111101100:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111101101:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111101110:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111101111:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111110000:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111110001:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111110010:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111110011:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111110100:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111110101:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111110110:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111110111:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111111000:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111111001:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111111010:	sigmoid_prime = 18'b000000000000011111;
		14'b10110111111011:	sigmoid_prime = 18'b000000000000100000;
		14'b10110111111100:	sigmoid_prime = 18'b000000000000100000;
		14'b10110111111101:	sigmoid_prime = 18'b000000000000100000;
		14'b10110111111110:	sigmoid_prime = 18'b000000000000100000;
		14'b10110111111111:	sigmoid_prime = 18'b000000000000100000;
		14'b10111000000000:	sigmoid_prime = 18'b000000000000100000;
		14'b10111000000001:	sigmoid_prime = 18'b000000000000100000;
		14'b10111000000010:	sigmoid_prime = 18'b000000000000100000;
		14'b10111000000011:	sigmoid_prime = 18'b000000000000100000;
		14'b10111000000100:	sigmoid_prime = 18'b000000000000100000;
		14'b10111000000101:	sigmoid_prime = 18'b000000000000100000;
		14'b10111000000110:	sigmoid_prime = 18'b000000000000100000;
		14'b10111000000111:	sigmoid_prime = 18'b000000000000100000;
		14'b10111000001000:	sigmoid_prime = 18'b000000000000100000;
		14'b10111000001001:	sigmoid_prime = 18'b000000000000100000;
		14'b10111000001010:	sigmoid_prime = 18'b000000000000100000;
		14'b10111000001011:	sigmoid_prime = 18'b000000000000100001;
		14'b10111000001100:	sigmoid_prime = 18'b000000000000100001;
		14'b10111000001101:	sigmoid_prime = 18'b000000000000100001;
		14'b10111000001110:	sigmoid_prime = 18'b000000000000100001;
		14'b10111000001111:	sigmoid_prime = 18'b000000000000100001;
		14'b10111000010000:	sigmoid_prime = 18'b000000000000100001;
		14'b10111000010001:	sigmoid_prime = 18'b000000000000100001;
		14'b10111000010010:	sigmoid_prime = 18'b000000000000100001;
		14'b10111000010011:	sigmoid_prime = 18'b000000000000100001;
		14'b10111000010100:	sigmoid_prime = 18'b000000000000100001;
		14'b10111000010101:	sigmoid_prime = 18'b000000000000100001;
		14'b10111000010110:	sigmoid_prime = 18'b000000000000100001;
		14'b10111000010111:	sigmoid_prime = 18'b000000000000100001;
		14'b10111000011000:	sigmoid_prime = 18'b000000000000100001;
		14'b10111000011001:	sigmoid_prime = 18'b000000000000100001;
		14'b10111000011010:	sigmoid_prime = 18'b000000000000100010;
		14'b10111000011011:	sigmoid_prime = 18'b000000000000100010;
		14'b10111000011100:	sigmoid_prime = 18'b000000000000100010;
		14'b10111000011101:	sigmoid_prime = 18'b000000000000100010;
		14'b10111000011110:	sigmoid_prime = 18'b000000000000100010;
		14'b10111000011111:	sigmoid_prime = 18'b000000000000100010;
		14'b10111000100000:	sigmoid_prime = 18'b000000000000100010;
		14'b10111000100001:	sigmoid_prime = 18'b000000000000100010;
		14'b10111000100010:	sigmoid_prime = 18'b000000000000100010;
		14'b10111000100011:	sigmoid_prime = 18'b000000000000100010;
		14'b10111000100100:	sigmoid_prime = 18'b000000000000100010;
		14'b10111000100101:	sigmoid_prime = 18'b000000000000100010;
		14'b10111000100110:	sigmoid_prime = 18'b000000000000100010;
		14'b10111000100111:	sigmoid_prime = 18'b000000000000100010;
		14'b10111000101000:	sigmoid_prime = 18'b000000000000100010;
		14'b10111000101001:	sigmoid_prime = 18'b000000000000100011;
		14'b10111000101010:	sigmoid_prime = 18'b000000000000100011;
		14'b10111000101011:	sigmoid_prime = 18'b000000000000100011;
		14'b10111000101100:	sigmoid_prime = 18'b000000000000100011;
		14'b10111000101101:	sigmoid_prime = 18'b000000000000100011;
		14'b10111000101110:	sigmoid_prime = 18'b000000000000100011;
		14'b10111000101111:	sigmoid_prime = 18'b000000000000100011;
		14'b10111000110000:	sigmoid_prime = 18'b000000000000100011;
		14'b10111000110001:	sigmoid_prime = 18'b000000000000100011;
		14'b10111000110010:	sigmoid_prime = 18'b000000000000100011;
		14'b10111000110011:	sigmoid_prime = 18'b000000000000100011;
		14'b10111000110100:	sigmoid_prime = 18'b000000000000100011;
		14'b10111000110101:	sigmoid_prime = 18'b000000000000100011;
		14'b10111000110110:	sigmoid_prime = 18'b000000000000100011;
		14'b10111000110111:	sigmoid_prime = 18'b000000000000100100;
		14'b10111000111000:	sigmoid_prime = 18'b000000000000100100;
		14'b10111000111001:	sigmoid_prime = 18'b000000000000100100;
		14'b10111000111010:	sigmoid_prime = 18'b000000000000100100;
		14'b10111000111011:	sigmoid_prime = 18'b000000000000100100;
		14'b10111000111100:	sigmoid_prime = 18'b000000000000100100;
		14'b10111000111101:	sigmoid_prime = 18'b000000000000100100;
		14'b10111000111110:	sigmoid_prime = 18'b000000000000100100;
		14'b10111000111111:	sigmoid_prime = 18'b000000000000100100;
		14'b10111001000000:	sigmoid_prime = 18'b000000000000100100;
		14'b10111001000001:	sigmoid_prime = 18'b000000000000100100;
		14'b10111001000010:	sigmoid_prime = 18'b000000000000100100;
		14'b10111001000011:	sigmoid_prime = 18'b000000000000100100;
		14'b10111001000100:	sigmoid_prime = 18'b000000000000100100;
		14'b10111001000101:	sigmoid_prime = 18'b000000000000100101;
		14'b10111001000110:	sigmoid_prime = 18'b000000000000100101;
		14'b10111001000111:	sigmoid_prime = 18'b000000000000100101;
		14'b10111001001000:	sigmoid_prime = 18'b000000000000100101;
		14'b10111001001001:	sigmoid_prime = 18'b000000000000100101;
		14'b10111001001010:	sigmoid_prime = 18'b000000000000100101;
		14'b10111001001011:	sigmoid_prime = 18'b000000000000100101;
		14'b10111001001100:	sigmoid_prime = 18'b000000000000100101;
		14'b10111001001101:	sigmoid_prime = 18'b000000000000100101;
		14'b10111001001110:	sigmoid_prime = 18'b000000000000100101;
		14'b10111001001111:	sigmoid_prime = 18'b000000000000100101;
		14'b10111001010000:	sigmoid_prime = 18'b000000000000100101;
		14'b10111001010001:	sigmoid_prime = 18'b000000000000100101;
		14'b10111001010010:	sigmoid_prime = 18'b000000000000100101;
		14'b10111001010011:	sigmoid_prime = 18'b000000000000100110;
		14'b10111001010100:	sigmoid_prime = 18'b000000000000100110;
		14'b10111001010101:	sigmoid_prime = 18'b000000000000100110;
		14'b10111001010110:	sigmoid_prime = 18'b000000000000100110;
		14'b10111001010111:	sigmoid_prime = 18'b000000000000100110;
		14'b10111001011000:	sigmoid_prime = 18'b000000000000100110;
		14'b10111001011001:	sigmoid_prime = 18'b000000000000100110;
		14'b10111001011010:	sigmoid_prime = 18'b000000000000100110;
		14'b10111001011011:	sigmoid_prime = 18'b000000000000100110;
		14'b10111001011100:	sigmoid_prime = 18'b000000000000100110;
		14'b10111001011101:	sigmoid_prime = 18'b000000000000100110;
		14'b10111001011110:	sigmoid_prime = 18'b000000000000100110;
		14'b10111001011111:	sigmoid_prime = 18'b000000000000100110;
		14'b10111001100000:	sigmoid_prime = 18'b000000000000100111;
		14'b10111001100001:	sigmoid_prime = 18'b000000000000100111;
		14'b10111001100010:	sigmoid_prime = 18'b000000000000100111;
		14'b10111001100011:	sigmoid_prime = 18'b000000000000100111;
		14'b10111001100100:	sigmoid_prime = 18'b000000000000100111;
		14'b10111001100101:	sigmoid_prime = 18'b000000000000100111;
		14'b10111001100110:	sigmoid_prime = 18'b000000000000100111;
		14'b10111001100111:	sigmoid_prime = 18'b000000000000100111;
		14'b10111001101000:	sigmoid_prime = 18'b000000000000100111;
		14'b10111001101001:	sigmoid_prime = 18'b000000000000100111;
		14'b10111001101010:	sigmoid_prime = 18'b000000000000100111;
		14'b10111001101011:	sigmoid_prime = 18'b000000000000100111;
		14'b10111001101100:	sigmoid_prime = 18'b000000000000100111;
		14'b10111001101101:	sigmoid_prime = 18'b000000000000101000;
		14'b10111001101110:	sigmoid_prime = 18'b000000000000101000;
		14'b10111001101111:	sigmoid_prime = 18'b000000000000101000;
		14'b10111001110000:	sigmoid_prime = 18'b000000000000101000;
		14'b10111001110001:	sigmoid_prime = 18'b000000000000101000;
		14'b10111001110010:	sigmoid_prime = 18'b000000000000101000;
		14'b10111001110011:	sigmoid_prime = 18'b000000000000101000;
		14'b10111001110100:	sigmoid_prime = 18'b000000000000101000;
		14'b10111001110101:	sigmoid_prime = 18'b000000000000101000;
		14'b10111001110110:	sigmoid_prime = 18'b000000000000101000;
		14'b10111001110111:	sigmoid_prime = 18'b000000000000101000;
		14'b10111001111000:	sigmoid_prime = 18'b000000000000101000;
		14'b10111001111001:	sigmoid_prime = 18'b000000000000101000;
		14'b10111001111010:	sigmoid_prime = 18'b000000000000101001;
		14'b10111001111011:	sigmoid_prime = 18'b000000000000101001;
		14'b10111001111100:	sigmoid_prime = 18'b000000000000101001;
		14'b10111001111101:	sigmoid_prime = 18'b000000000000101001;
		14'b10111001111110:	sigmoid_prime = 18'b000000000000101001;
		14'b10111001111111:	sigmoid_prime = 18'b000000000000101001;
		14'b10111010000000:	sigmoid_prime = 18'b000000000000101001;
		14'b10111010000001:	sigmoid_prime = 18'b000000000000101001;
		14'b10111010000010:	sigmoid_prime = 18'b000000000000101001;
		14'b10111010000011:	sigmoid_prime = 18'b000000000000101001;
		14'b10111010000100:	sigmoid_prime = 18'b000000000000101001;
		14'b10111010000101:	sigmoid_prime = 18'b000000000000101001;
		14'b10111010000110:	sigmoid_prime = 18'b000000000000101010;
		14'b10111010000111:	sigmoid_prime = 18'b000000000000101010;
		14'b10111010001000:	sigmoid_prime = 18'b000000000000101010;
		14'b10111010001001:	sigmoid_prime = 18'b000000000000101010;
		14'b10111010001010:	sigmoid_prime = 18'b000000000000101010;
		14'b10111010001011:	sigmoid_prime = 18'b000000000000101010;
		14'b10111010001100:	sigmoid_prime = 18'b000000000000101010;
		14'b10111010001101:	sigmoid_prime = 18'b000000000000101010;
		14'b10111010001110:	sigmoid_prime = 18'b000000000000101010;
		14'b10111010001111:	sigmoid_prime = 18'b000000000000101010;
		14'b10111010010000:	sigmoid_prime = 18'b000000000000101010;
		14'b10111010010001:	sigmoid_prime = 18'b000000000000101010;
		14'b10111010010010:	sigmoid_prime = 18'b000000000000101011;
		14'b10111010010011:	sigmoid_prime = 18'b000000000000101011;
		14'b10111010010100:	sigmoid_prime = 18'b000000000000101011;
		14'b10111010010101:	sigmoid_prime = 18'b000000000000101011;
		14'b10111010010110:	sigmoid_prime = 18'b000000000000101011;
		14'b10111010010111:	sigmoid_prime = 18'b000000000000101011;
		14'b10111010011000:	sigmoid_prime = 18'b000000000000101011;
		14'b10111010011001:	sigmoid_prime = 18'b000000000000101011;
		14'b10111010011010:	sigmoid_prime = 18'b000000000000101011;
		14'b10111010011011:	sigmoid_prime = 18'b000000000000101011;
		14'b10111010011100:	sigmoid_prime = 18'b000000000000101011;
		14'b10111010011101:	sigmoid_prime = 18'b000000000000101011;
		14'b10111010011110:	sigmoid_prime = 18'b000000000000101100;
		14'b10111010011111:	sigmoid_prime = 18'b000000000000101100;
		14'b10111010100000:	sigmoid_prime = 18'b000000000000101100;
		14'b10111010100001:	sigmoid_prime = 18'b000000000000101100;
		14'b10111010100010:	sigmoid_prime = 18'b000000000000101100;
		14'b10111010100011:	sigmoid_prime = 18'b000000000000101100;
		14'b10111010100100:	sigmoid_prime = 18'b000000000000101100;
		14'b10111010100101:	sigmoid_prime = 18'b000000000000101100;
		14'b10111010100110:	sigmoid_prime = 18'b000000000000101100;
		14'b10111010100111:	sigmoid_prime = 18'b000000000000101100;
		14'b10111010101000:	sigmoid_prime = 18'b000000000000101100;
		14'b10111010101001:	sigmoid_prime = 18'b000000000000101100;
		14'b10111010101010:	sigmoid_prime = 18'b000000000000101101;
		14'b10111010101011:	sigmoid_prime = 18'b000000000000101101;
		14'b10111010101100:	sigmoid_prime = 18'b000000000000101101;
		14'b10111010101101:	sigmoid_prime = 18'b000000000000101101;
		14'b10111010101110:	sigmoid_prime = 18'b000000000000101101;
		14'b10111010101111:	sigmoid_prime = 18'b000000000000101101;
		14'b10111010110000:	sigmoid_prime = 18'b000000000000101101;
		14'b10111010110001:	sigmoid_prime = 18'b000000000000101101;
		14'b10111010110010:	sigmoid_prime = 18'b000000000000101101;
		14'b10111010110011:	sigmoid_prime = 18'b000000000000101101;
		14'b10111010110100:	sigmoid_prime = 18'b000000000000101101;
		14'b10111010110101:	sigmoid_prime = 18'b000000000000101110;
		14'b10111010110110:	sigmoid_prime = 18'b000000000000101110;
		14'b10111010110111:	sigmoid_prime = 18'b000000000000101110;
		14'b10111010111000:	sigmoid_prime = 18'b000000000000101110;
		14'b10111010111001:	sigmoid_prime = 18'b000000000000101110;
		14'b10111010111010:	sigmoid_prime = 18'b000000000000101110;
		14'b10111010111011:	sigmoid_prime = 18'b000000000000101110;
		14'b10111010111100:	sigmoid_prime = 18'b000000000000101110;
		14'b10111010111101:	sigmoid_prime = 18'b000000000000101110;
		14'b10111010111110:	sigmoid_prime = 18'b000000000000101110;
		14'b10111010111111:	sigmoid_prime = 18'b000000000000101110;
		14'b10111011000000:	sigmoid_prime = 18'b000000000000101111;
		14'b10111011000001:	sigmoid_prime = 18'b000000000000101111;
		14'b10111011000010:	sigmoid_prime = 18'b000000000000101111;
		14'b10111011000011:	sigmoid_prime = 18'b000000000000101111;
		14'b10111011000100:	sigmoid_prime = 18'b000000000000101111;
		14'b10111011000101:	sigmoid_prime = 18'b000000000000101111;
		14'b10111011000110:	sigmoid_prime = 18'b000000000000101111;
		14'b10111011000111:	sigmoid_prime = 18'b000000000000101111;
		14'b10111011001000:	sigmoid_prime = 18'b000000000000101111;
		14'b10111011001001:	sigmoid_prime = 18'b000000000000101111;
		14'b10111011001010:	sigmoid_prime = 18'b000000000000101111;
		14'b10111011001011:	sigmoid_prime = 18'b000000000000110000;
		14'b10111011001100:	sigmoid_prime = 18'b000000000000110000;
		14'b10111011001101:	sigmoid_prime = 18'b000000000000110000;
		14'b10111011001110:	sigmoid_prime = 18'b000000000000110000;
		14'b10111011001111:	sigmoid_prime = 18'b000000000000110000;
		14'b10111011010000:	sigmoid_prime = 18'b000000000000110000;
		14'b10111011010001:	sigmoid_prime = 18'b000000000000110000;
		14'b10111011010010:	sigmoid_prime = 18'b000000000000110000;
		14'b10111011010011:	sigmoid_prime = 18'b000000000000110000;
		14'b10111011010100:	sigmoid_prime = 18'b000000000000110000;
		14'b10111011010101:	sigmoid_prime = 18'b000000000000110001;
		14'b10111011010110:	sigmoid_prime = 18'b000000000000110001;
		14'b10111011010111:	sigmoid_prime = 18'b000000000000110001;
		14'b10111011011000:	sigmoid_prime = 18'b000000000000110001;
		14'b10111011011001:	sigmoid_prime = 18'b000000000000110001;
		14'b10111011011010:	sigmoid_prime = 18'b000000000000110001;
		14'b10111011011011:	sigmoid_prime = 18'b000000000000110001;
		14'b10111011011100:	sigmoid_prime = 18'b000000000000110001;
		14'b10111011011101:	sigmoid_prime = 18'b000000000000110001;
		14'b10111011011110:	sigmoid_prime = 18'b000000000000110001;
		14'b10111011011111:	sigmoid_prime = 18'b000000000000110001;
		14'b10111011100000:	sigmoid_prime = 18'b000000000000110010;
		14'b10111011100001:	sigmoid_prime = 18'b000000000000110010;
		14'b10111011100010:	sigmoid_prime = 18'b000000000000110010;
		14'b10111011100011:	sigmoid_prime = 18'b000000000000110010;
		14'b10111011100100:	sigmoid_prime = 18'b000000000000110010;
		14'b10111011100101:	sigmoid_prime = 18'b000000000000110010;
		14'b10111011100110:	sigmoid_prime = 18'b000000000000110010;
		14'b10111011100111:	sigmoid_prime = 18'b000000000000110010;
		14'b10111011101000:	sigmoid_prime = 18'b000000000000110010;
		14'b10111011101001:	sigmoid_prime = 18'b000000000000110010;
		14'b10111011101010:	sigmoid_prime = 18'b000000000000110011;
		14'b10111011101011:	sigmoid_prime = 18'b000000000000110011;
		14'b10111011101100:	sigmoid_prime = 18'b000000000000110011;
		14'b10111011101101:	sigmoid_prime = 18'b000000000000110011;
		14'b10111011101110:	sigmoid_prime = 18'b000000000000110011;
		14'b10111011101111:	sigmoid_prime = 18'b000000000000110011;
		14'b10111011110000:	sigmoid_prime = 18'b000000000000110011;
		14'b10111011110001:	sigmoid_prime = 18'b000000000000110011;
		14'b10111011110010:	sigmoid_prime = 18'b000000000000110011;
		14'b10111011110011:	sigmoid_prime = 18'b000000000000110011;
		14'b10111011110100:	sigmoid_prime = 18'b000000000000110100;
		14'b10111011110101:	sigmoid_prime = 18'b000000000000110100;
		14'b10111011110110:	sigmoid_prime = 18'b000000000000110100;
		14'b10111011110111:	sigmoid_prime = 18'b000000000000110100;
		14'b10111011111000:	sigmoid_prime = 18'b000000000000110100;
		14'b10111011111001:	sigmoid_prime = 18'b000000000000110100;
		14'b10111011111010:	sigmoid_prime = 18'b000000000000110100;
		14'b10111011111011:	sigmoid_prime = 18'b000000000000110100;
		14'b10111011111100:	sigmoid_prime = 18'b000000000000110100;
		14'b10111011111101:	sigmoid_prime = 18'b000000000000110101;
		14'b10111011111110:	sigmoid_prime = 18'b000000000000110101;
		14'b10111011111111:	sigmoid_prime = 18'b000000000000110101;
		14'b10111100000000:	sigmoid_prime = 18'b000000000000110101;
		14'b10111100000001:	sigmoid_prime = 18'b000000000000110101;
		14'b10111100000010:	sigmoid_prime = 18'b000000000000110101;
		14'b10111100000011:	sigmoid_prime = 18'b000000000000110101;
		14'b10111100000100:	sigmoid_prime = 18'b000000000000110101;
		14'b10111100000101:	sigmoid_prime = 18'b000000000000110101;
		14'b10111100000110:	sigmoid_prime = 18'b000000000000110101;
		14'b10111100000111:	sigmoid_prime = 18'b000000000000110110;
		14'b10111100001000:	sigmoid_prime = 18'b000000000000110110;
		14'b10111100001001:	sigmoid_prime = 18'b000000000000110110;
		14'b10111100001010:	sigmoid_prime = 18'b000000000000110110;
		14'b10111100001011:	sigmoid_prime = 18'b000000000000110110;
		14'b10111100001100:	sigmoid_prime = 18'b000000000000110110;
		14'b10111100001101:	sigmoid_prime = 18'b000000000000110110;
		14'b10111100001110:	sigmoid_prime = 18'b000000000000110110;
		14'b10111100001111:	sigmoid_prime = 18'b000000000000110110;
		14'b10111100010000:	sigmoid_prime = 18'b000000000000110111;
		14'b10111100010001:	sigmoid_prime = 18'b000000000000110111;
		14'b10111100010010:	sigmoid_prime = 18'b000000000000110111;
		14'b10111100010011:	sigmoid_prime = 18'b000000000000110111;
		14'b10111100010100:	sigmoid_prime = 18'b000000000000110111;
		14'b10111100010101:	sigmoid_prime = 18'b000000000000110111;
		14'b10111100010110:	sigmoid_prime = 18'b000000000000110111;
		14'b10111100010111:	sigmoid_prime = 18'b000000000000110111;
		14'b10111100011000:	sigmoid_prime = 18'b000000000000110111;
		14'b10111100011001:	sigmoid_prime = 18'b000000000000110111;
		14'b10111100011010:	sigmoid_prime = 18'b000000000000111000;
		14'b10111100011011:	sigmoid_prime = 18'b000000000000111000;
		14'b10111100011100:	sigmoid_prime = 18'b000000000000111000;
		14'b10111100011101:	sigmoid_prime = 18'b000000000000111000;
		14'b10111100011110:	sigmoid_prime = 18'b000000000000111000;
		14'b10111100011111:	sigmoid_prime = 18'b000000000000111000;
		14'b10111100100000:	sigmoid_prime = 18'b000000000000111000;
		14'b10111100100001:	sigmoid_prime = 18'b000000000000111000;
		14'b10111100100010:	sigmoid_prime = 18'b000000000000111000;
		14'b10111100100011:	sigmoid_prime = 18'b000000000000111001;
		14'b10111100100100:	sigmoid_prime = 18'b000000000000111001;
		14'b10111100100101:	sigmoid_prime = 18'b000000000000111001;
		14'b10111100100110:	sigmoid_prime = 18'b000000000000111001;
		14'b10111100100111:	sigmoid_prime = 18'b000000000000111001;
		14'b10111100101000:	sigmoid_prime = 18'b000000000000111001;
		14'b10111100101001:	sigmoid_prime = 18'b000000000000111001;
		14'b10111100101010:	sigmoid_prime = 18'b000000000000111001;
		14'b10111100101011:	sigmoid_prime = 18'b000000000000111001;
		14'b10111100101100:	sigmoid_prime = 18'b000000000000111010;
		14'b10111100101101:	sigmoid_prime = 18'b000000000000111010;
		14'b10111100101110:	sigmoid_prime = 18'b000000000000111010;
		14'b10111100101111:	sigmoid_prime = 18'b000000000000111010;
		14'b10111100110000:	sigmoid_prime = 18'b000000000000111010;
		14'b10111100110001:	sigmoid_prime = 18'b000000000000111010;
		14'b10111100110010:	sigmoid_prime = 18'b000000000000111010;
		14'b10111100110011:	sigmoid_prime = 18'b000000000000111010;
		14'b10111100110100:	sigmoid_prime = 18'b000000000000111011;
		14'b10111100110101:	sigmoid_prime = 18'b000000000000111011;
		14'b10111100110110:	sigmoid_prime = 18'b000000000000111011;
		14'b10111100110111:	sigmoid_prime = 18'b000000000000111011;
		14'b10111100111000:	sigmoid_prime = 18'b000000000000111011;
		14'b10111100111001:	sigmoid_prime = 18'b000000000000111011;
		14'b10111100111010:	sigmoid_prime = 18'b000000000000111011;
		14'b10111100111011:	sigmoid_prime = 18'b000000000000111011;
		14'b10111100111100:	sigmoid_prime = 18'b000000000000111011;
		14'b10111100111101:	sigmoid_prime = 18'b000000000000111100;
		14'b10111100111110:	sigmoid_prime = 18'b000000000000111100;
		14'b10111100111111:	sigmoid_prime = 18'b000000000000111100;
		14'b10111101000000:	sigmoid_prime = 18'b000000000000111100;
		14'b10111101000001:	sigmoid_prime = 18'b000000000000111100;
		14'b10111101000010:	sigmoid_prime = 18'b000000000000111100;
		14'b10111101000011:	sigmoid_prime = 18'b000000000000111100;
		14'b10111101000100:	sigmoid_prime = 18'b000000000000111100;
		14'b10111101000101:	sigmoid_prime = 18'b000000000000111101;
		14'b10111101000110:	sigmoid_prime = 18'b000000000000111101;
		14'b10111101000111:	sigmoid_prime = 18'b000000000000111101;
		14'b10111101001000:	sigmoid_prime = 18'b000000000000111101;
		14'b10111101001001:	sigmoid_prime = 18'b000000000000111101;
		14'b10111101001010:	sigmoid_prime = 18'b000000000000111101;
		14'b10111101001011:	sigmoid_prime = 18'b000000000000111101;
		14'b10111101001100:	sigmoid_prime = 18'b000000000000111101;
		14'b10111101001101:	sigmoid_prime = 18'b000000000000111101;
		14'b10111101001110:	sigmoid_prime = 18'b000000000000111110;
		14'b10111101001111:	sigmoid_prime = 18'b000000000000111110;
		14'b10111101010000:	sigmoid_prime = 18'b000000000000111110;
		14'b10111101010001:	sigmoid_prime = 18'b000000000000111110;
		14'b10111101010010:	sigmoid_prime = 18'b000000000000111110;
		14'b10111101010011:	sigmoid_prime = 18'b000000000000111110;
		14'b10111101010100:	sigmoid_prime = 18'b000000000000111110;
		14'b10111101010101:	sigmoid_prime = 18'b000000000000111110;
		14'b10111101010110:	sigmoid_prime = 18'b000000000000111111;
		14'b10111101010111:	sigmoid_prime = 18'b000000000000111111;
		14'b10111101011000:	sigmoid_prime = 18'b000000000000111111;
		14'b10111101011001:	sigmoid_prime = 18'b000000000000111111;
		14'b10111101011010:	sigmoid_prime = 18'b000000000000111111;
		14'b10111101011011:	sigmoid_prime = 18'b000000000000111111;
		14'b10111101011100:	sigmoid_prime = 18'b000000000000111111;
		14'b10111101011101:	sigmoid_prime = 18'b000000000000111111;
		14'b10111101011110:	sigmoid_prime = 18'b000000000001000000;
		14'b10111101011111:	sigmoid_prime = 18'b000000000001000000;
		14'b10111101100000:	sigmoid_prime = 18'b000000000001000000;
		14'b10111101100001:	sigmoid_prime = 18'b000000000001000000;
		14'b10111101100010:	sigmoid_prime = 18'b000000000001000000;
		14'b10111101100011:	sigmoid_prime = 18'b000000000001000000;
		14'b10111101100100:	sigmoid_prime = 18'b000000000001000000;
		14'b10111101100101:	sigmoid_prime = 18'b000000000001000000;
		14'b10111101100110:	sigmoid_prime = 18'b000000000001000001;
		14'b10111101100111:	sigmoid_prime = 18'b000000000001000001;
		14'b10111101101000:	sigmoid_prime = 18'b000000000001000001;
		14'b10111101101001:	sigmoid_prime = 18'b000000000001000001;
		14'b10111101101010:	sigmoid_prime = 18'b000000000001000001;
		14'b10111101101011:	sigmoid_prime = 18'b000000000001000001;
		14'b10111101101100:	sigmoid_prime = 18'b000000000001000001;
		14'b10111101101101:	sigmoid_prime = 18'b000000000001000001;
		14'b10111101101110:	sigmoid_prime = 18'b000000000001000010;
		14'b10111101101111:	sigmoid_prime = 18'b000000000001000010;
		14'b10111101110000:	sigmoid_prime = 18'b000000000001000010;
		14'b10111101110001:	sigmoid_prime = 18'b000000000001000010;
		14'b10111101110010:	sigmoid_prime = 18'b000000000001000010;
		14'b10111101110011:	sigmoid_prime = 18'b000000000001000010;
		14'b10111101110100:	sigmoid_prime = 18'b000000000001000010;
		14'b10111101110101:	sigmoid_prime = 18'b000000000001000010;
		14'b10111101110110:	sigmoid_prime = 18'b000000000001000011;
		14'b10111101110111:	sigmoid_prime = 18'b000000000001000011;
		14'b10111101111000:	sigmoid_prime = 18'b000000000001000011;
		14'b10111101111001:	sigmoid_prime = 18'b000000000001000011;
		14'b10111101111010:	sigmoid_prime = 18'b000000000001000011;
		14'b10111101111011:	sigmoid_prime = 18'b000000000001000011;
		14'b10111101111100:	sigmoid_prime = 18'b000000000001000011;
		14'b10111101111101:	sigmoid_prime = 18'b000000000001000100;
		14'b10111101111110:	sigmoid_prime = 18'b000000000001000100;
		14'b10111101111111:	sigmoid_prime = 18'b000000000001000100;
		14'b10111110000000:	sigmoid_prime = 18'b000000000001000100;
		14'b10111110000001:	sigmoid_prime = 18'b000000000001000100;
		14'b10111110000010:	sigmoid_prime = 18'b000000000001000100;
		14'b10111110000011:	sigmoid_prime = 18'b000000000001000100;
		14'b10111110000100:	sigmoid_prime = 18'b000000000001000100;
		14'b10111110000101:	sigmoid_prime = 18'b000000000001000101;
		14'b10111110000110:	sigmoid_prime = 18'b000000000001000101;
		14'b10111110000111:	sigmoid_prime = 18'b000000000001000101;
		14'b10111110001000:	sigmoid_prime = 18'b000000000001000101;
		14'b10111110001001:	sigmoid_prime = 18'b000000000001000101;
		14'b10111110001010:	sigmoid_prime = 18'b000000000001000101;
		14'b10111110001011:	sigmoid_prime = 18'b000000000001000101;
		14'b10111110001100:	sigmoid_prime = 18'b000000000001000110;
		14'b10111110001101:	sigmoid_prime = 18'b000000000001000110;
		14'b10111110001110:	sigmoid_prime = 18'b000000000001000110;
		14'b10111110001111:	sigmoid_prime = 18'b000000000001000110;
		14'b10111110010000:	sigmoid_prime = 18'b000000000001000110;
		14'b10111110010001:	sigmoid_prime = 18'b000000000001000110;
		14'b10111110010010:	sigmoid_prime = 18'b000000000001000110;
		14'b10111110010011:	sigmoid_prime = 18'b000000000001000111;
		14'b10111110010100:	sigmoid_prime = 18'b000000000001000111;
		14'b10111110010101:	sigmoid_prime = 18'b000000000001000111;
		14'b10111110010110:	sigmoid_prime = 18'b000000000001000111;
		14'b10111110010111:	sigmoid_prime = 18'b000000000001000111;
		14'b10111110011000:	sigmoid_prime = 18'b000000000001000111;
		14'b10111110011001:	sigmoid_prime = 18'b000000000001000111;
		14'b10111110011010:	sigmoid_prime = 18'b000000000001001000;
		14'b10111110011011:	sigmoid_prime = 18'b000000000001001000;
		14'b10111110011100:	sigmoid_prime = 18'b000000000001001000;
		14'b10111110011101:	sigmoid_prime = 18'b000000000001001000;
		14'b10111110011110:	sigmoid_prime = 18'b000000000001001000;
		14'b10111110011111:	sigmoid_prime = 18'b000000000001001000;
		14'b10111110100000:	sigmoid_prime = 18'b000000000001001000;
		14'b10111110100001:	sigmoid_prime = 18'b000000000001001001;
		14'b10111110100010:	sigmoid_prime = 18'b000000000001001001;
		14'b10111110100011:	sigmoid_prime = 18'b000000000001001001;
		14'b10111110100100:	sigmoid_prime = 18'b000000000001001001;
		14'b10111110100101:	sigmoid_prime = 18'b000000000001001001;
		14'b10111110100110:	sigmoid_prime = 18'b000000000001001001;
		14'b10111110100111:	sigmoid_prime = 18'b000000000001001001;
		14'b10111110101000:	sigmoid_prime = 18'b000000000001001010;
		14'b10111110101001:	sigmoid_prime = 18'b000000000001001010;
		14'b10111110101010:	sigmoid_prime = 18'b000000000001001010;
		14'b10111110101011:	sigmoid_prime = 18'b000000000001001010;
		14'b10111110101100:	sigmoid_prime = 18'b000000000001001010;
		14'b10111110101101:	sigmoid_prime = 18'b000000000001001010;
		14'b10111110101110:	sigmoid_prime = 18'b000000000001001010;
		14'b10111110101111:	sigmoid_prime = 18'b000000000001001011;
		14'b10111110110000:	sigmoid_prime = 18'b000000000001001011;
		14'b10111110110001:	sigmoid_prime = 18'b000000000001001011;
		14'b10111110110010:	sigmoid_prime = 18'b000000000001001011;
		14'b10111110110011:	sigmoid_prime = 18'b000000000001001011;
		14'b10111110110100:	sigmoid_prime = 18'b000000000001001011;
		14'b10111110110101:	sigmoid_prime = 18'b000000000001001011;
		14'b10111110110110:	sigmoid_prime = 18'b000000000001001100;
		14'b10111110110111:	sigmoid_prime = 18'b000000000001001100;
		14'b10111110111000:	sigmoid_prime = 18'b000000000001001100;
		14'b10111110111001:	sigmoid_prime = 18'b000000000001001100;
		14'b10111110111010:	sigmoid_prime = 18'b000000000001001100;
		14'b10111110111011:	sigmoid_prime = 18'b000000000001001100;
		14'b10111110111100:	sigmoid_prime = 18'b000000000001001100;
		14'b10111110111101:	sigmoid_prime = 18'b000000000001001101;
		14'b10111110111110:	sigmoid_prime = 18'b000000000001001101;
		14'b10111110111111:	sigmoid_prime = 18'b000000000001001101;
		14'b10111111000000:	sigmoid_prime = 18'b000000000001001101;
		14'b10111111000001:	sigmoid_prime = 18'b000000000001001101;
		14'b10111111000010:	sigmoid_prime = 18'b000000000001001101;
		14'b10111111000011:	sigmoid_prime = 18'b000000000001001110;
		14'b10111111000100:	sigmoid_prime = 18'b000000000001001110;
		14'b10111111000101:	sigmoid_prime = 18'b000000000001001110;
		14'b10111111000110:	sigmoid_prime = 18'b000000000001001110;
		14'b10111111000111:	sigmoid_prime = 18'b000000000001001110;
		14'b10111111001000:	sigmoid_prime = 18'b000000000001001110;
		14'b10111111001001:	sigmoid_prime = 18'b000000000001001110;
		14'b10111111001010:	sigmoid_prime = 18'b000000000001001111;
		14'b10111111001011:	sigmoid_prime = 18'b000000000001001111;
		14'b10111111001100:	sigmoid_prime = 18'b000000000001001111;
		14'b10111111001101:	sigmoid_prime = 18'b000000000001001111;
		14'b10111111001110:	sigmoid_prime = 18'b000000000001001111;
		14'b10111111001111:	sigmoid_prime = 18'b000000000001001111;
		14'b10111111010000:	sigmoid_prime = 18'b000000000001010000;
		14'b10111111010001:	sigmoid_prime = 18'b000000000001010000;
		14'b10111111010010:	sigmoid_prime = 18'b000000000001010000;
		14'b10111111010011:	sigmoid_prime = 18'b000000000001010000;
		14'b10111111010100:	sigmoid_prime = 18'b000000000001010000;
		14'b10111111010101:	sigmoid_prime = 18'b000000000001010000;
		14'b10111111010110:	sigmoid_prime = 18'b000000000001010000;
		14'b10111111010111:	sigmoid_prime = 18'b000000000001010001;
		14'b10111111011000:	sigmoid_prime = 18'b000000000001010001;
		14'b10111111011001:	sigmoid_prime = 18'b000000000001010001;
		14'b10111111011010:	sigmoid_prime = 18'b000000000001010001;
		14'b10111111011011:	sigmoid_prime = 18'b000000000001010001;
		14'b10111111011100:	sigmoid_prime = 18'b000000000001010001;
		14'b10111111011101:	sigmoid_prime = 18'b000000000001010010;
		14'b10111111011110:	sigmoid_prime = 18'b000000000001010010;
		14'b10111111011111:	sigmoid_prime = 18'b000000000001010010;
		14'b10111111100000:	sigmoid_prime = 18'b000000000001010010;
		14'b10111111100001:	sigmoid_prime = 18'b000000000001010010;
		14'b10111111100010:	sigmoid_prime = 18'b000000000001010010;
		14'b10111111100011:	sigmoid_prime = 18'b000000000001010011;
		14'b10111111100100:	sigmoid_prime = 18'b000000000001010011;
		14'b10111111100101:	sigmoid_prime = 18'b000000000001010011;
		14'b10111111100110:	sigmoid_prime = 18'b000000000001010011;
		14'b10111111100111:	sigmoid_prime = 18'b000000000001010011;
		14'b10111111101000:	sigmoid_prime = 18'b000000000001010011;
		14'b10111111101001:	sigmoid_prime = 18'b000000000001010100;
		14'b10111111101010:	sigmoid_prime = 18'b000000000001010100;
		14'b10111111101011:	sigmoid_prime = 18'b000000000001010100;
		14'b10111111101100:	sigmoid_prime = 18'b000000000001010100;
		14'b10111111101101:	sigmoid_prime = 18'b000000000001010100;
		14'b10111111101110:	sigmoid_prime = 18'b000000000001010100;
		14'b10111111101111:	sigmoid_prime = 18'b000000000001010101;
		14'b10111111110000:	sigmoid_prime = 18'b000000000001010101;
		14'b10111111110001:	sigmoid_prime = 18'b000000000001010101;
		14'b10111111110010:	sigmoid_prime = 18'b000000000001010101;
		14'b10111111110011:	sigmoid_prime = 18'b000000000001010101;
		14'b10111111110100:	sigmoid_prime = 18'b000000000001010101;
		14'b10111111110101:	sigmoid_prime = 18'b000000000001010110;
		14'b10111111110110:	sigmoid_prime = 18'b000000000001010110;
		14'b10111111110111:	sigmoid_prime = 18'b000000000001010110;
		14'b10111111111000:	sigmoid_prime = 18'b000000000001010110;
		14'b10111111111001:	sigmoid_prime = 18'b000000000001010110;
		14'b10111111111010:	sigmoid_prime = 18'b000000000001010110;
		14'b10111111111011:	sigmoid_prime = 18'b000000000001010111;
		14'b10111111111100:	sigmoid_prime = 18'b000000000001010111;
		14'b10111111111101:	sigmoid_prime = 18'b000000000001010111;
		14'b10111111111110:	sigmoid_prime = 18'b000000000001010111;
		14'b10111111111111:	sigmoid_prime = 18'b000000000001010111;
		14'b11000000000000:	sigmoid_prime = 18'b000000000001010111;
		14'b11000000000001:	sigmoid_prime = 18'b000000000001011000;
		14'b11000000000010:	sigmoid_prime = 18'b000000000001011000;
		14'b11000000000011:	sigmoid_prime = 18'b000000000001011000;
		14'b11000000000100:	sigmoid_prime = 18'b000000000001011000;
		14'b11000000000101:	sigmoid_prime = 18'b000000000001011000;
		14'b11000000000110:	sigmoid_prime = 18'b000000000001011000;
		14'b11000000000111:	sigmoid_prime = 18'b000000000001011001;
		14'b11000000001000:	sigmoid_prime = 18'b000000000001011001;
		14'b11000000001001:	sigmoid_prime = 18'b000000000001011001;
		14'b11000000001010:	sigmoid_prime = 18'b000000000001011001;
		14'b11000000001011:	sigmoid_prime = 18'b000000000001011001;
		14'b11000000001100:	sigmoid_prime = 18'b000000000001011001;
		14'b11000000001101:	sigmoid_prime = 18'b000000000001011010;
		14'b11000000001110:	sigmoid_prime = 18'b000000000001011010;
		14'b11000000001111:	sigmoid_prime = 18'b000000000001011010;
		14'b11000000010000:	sigmoid_prime = 18'b000000000001011010;
		14'b11000000010001:	sigmoid_prime = 18'b000000000001011010;
		14'b11000000010010:	sigmoid_prime = 18'b000000000001011011;
		14'b11000000010011:	sigmoid_prime = 18'b000000000001011011;
		14'b11000000010100:	sigmoid_prime = 18'b000000000001011011;
		14'b11000000010101:	sigmoid_prime = 18'b000000000001011011;
		14'b11000000010110:	sigmoid_prime = 18'b000000000001011011;
		14'b11000000010111:	sigmoid_prime = 18'b000000000001011011;
		14'b11000000011000:	sigmoid_prime = 18'b000000000001011100;
		14'b11000000011001:	sigmoid_prime = 18'b000000000001011100;
		14'b11000000011010:	sigmoid_prime = 18'b000000000001011100;
		14'b11000000011011:	sigmoid_prime = 18'b000000000001011100;
		14'b11000000011100:	sigmoid_prime = 18'b000000000001011100;
		14'b11000000011101:	sigmoid_prime = 18'b000000000001011100;
		14'b11000000011110:	sigmoid_prime = 18'b000000000001011101;
		14'b11000000011111:	sigmoid_prime = 18'b000000000001011101;
		14'b11000000100000:	sigmoid_prime = 18'b000000000001011101;
		14'b11000000100001:	sigmoid_prime = 18'b000000000001011101;
		14'b11000000100010:	sigmoid_prime = 18'b000000000001011101;
		14'b11000000100011:	sigmoid_prime = 18'b000000000001011110;
		14'b11000000100100:	sigmoid_prime = 18'b000000000001011110;
		14'b11000000100101:	sigmoid_prime = 18'b000000000001011110;
		14'b11000000100110:	sigmoid_prime = 18'b000000000001011110;
		14'b11000000100111:	sigmoid_prime = 18'b000000000001011110;
		14'b11000000101000:	sigmoid_prime = 18'b000000000001011111;
		14'b11000000101001:	sigmoid_prime = 18'b000000000001011111;
		14'b11000000101010:	sigmoid_prime = 18'b000000000001011111;
		14'b11000000101011:	sigmoid_prime = 18'b000000000001011111;
		14'b11000000101100:	sigmoid_prime = 18'b000000000001011111;
		14'b11000000101101:	sigmoid_prime = 18'b000000000001011111;
		14'b11000000101110:	sigmoid_prime = 18'b000000000001100000;
		14'b11000000101111:	sigmoid_prime = 18'b000000000001100000;
		14'b11000000110000:	sigmoid_prime = 18'b000000000001100000;
		14'b11000000110001:	sigmoid_prime = 18'b000000000001100000;
		14'b11000000110010:	sigmoid_prime = 18'b000000000001100000;
		14'b11000000110011:	sigmoid_prime = 18'b000000000001100001;
		14'b11000000110100:	sigmoid_prime = 18'b000000000001100001;
		14'b11000000110101:	sigmoid_prime = 18'b000000000001100001;
		14'b11000000110110:	sigmoid_prime = 18'b000000000001100001;
		14'b11000000110111:	sigmoid_prime = 18'b000000000001100001;
		14'b11000000111000:	sigmoid_prime = 18'b000000000001100010;
		14'b11000000111001:	sigmoid_prime = 18'b000000000001100010;
		14'b11000000111010:	sigmoid_prime = 18'b000000000001100010;
		14'b11000000111011:	sigmoid_prime = 18'b000000000001100010;
		14'b11000000111100:	sigmoid_prime = 18'b000000000001100010;
		14'b11000000111101:	sigmoid_prime = 18'b000000000001100010;
		14'b11000000111110:	sigmoid_prime = 18'b000000000001100011;
		14'b11000000111111:	sigmoid_prime = 18'b000000000001100011;
		14'b11000001000000:	sigmoid_prime = 18'b000000000001100011;
		14'b11000001000001:	sigmoid_prime = 18'b000000000001100011;
		14'b11000001000010:	sigmoid_prime = 18'b000000000001100011;
		14'b11000001000011:	sigmoid_prime = 18'b000000000001100100;
		14'b11000001000100:	sigmoid_prime = 18'b000000000001100100;
		14'b11000001000101:	sigmoid_prime = 18'b000000000001100100;
		14'b11000001000110:	sigmoid_prime = 18'b000000000001100100;
		14'b11000001000111:	sigmoid_prime = 18'b000000000001100100;
		14'b11000001001000:	sigmoid_prime = 18'b000000000001100101;
		14'b11000001001001:	sigmoid_prime = 18'b000000000001100101;
		14'b11000001001010:	sigmoid_prime = 18'b000000000001100101;
		14'b11000001001011:	sigmoid_prime = 18'b000000000001100101;
		14'b11000001001100:	sigmoid_prime = 18'b000000000001100101;
		14'b11000001001101:	sigmoid_prime = 18'b000000000001100110;
		14'b11000001001110:	sigmoid_prime = 18'b000000000001100110;
		14'b11000001001111:	sigmoid_prime = 18'b000000000001100110;
		14'b11000001010000:	sigmoid_prime = 18'b000000000001100110;
		14'b11000001010001:	sigmoid_prime = 18'b000000000001100110;
		14'b11000001010010:	sigmoid_prime = 18'b000000000001100111;
		14'b11000001010011:	sigmoid_prime = 18'b000000000001100111;
		14'b11000001010100:	sigmoid_prime = 18'b000000000001100111;
		14'b11000001010101:	sigmoid_prime = 18'b000000000001100111;
		14'b11000001010110:	sigmoid_prime = 18'b000000000001100111;
		14'b11000001010111:	sigmoid_prime = 18'b000000000001101000;
		14'b11000001011000:	sigmoid_prime = 18'b000000000001101000;
		14'b11000001011001:	sigmoid_prime = 18'b000000000001101000;
		14'b11000001011010:	sigmoid_prime = 18'b000000000001101000;
		14'b11000001011011:	sigmoid_prime = 18'b000000000001101000;
		14'b11000001011100:	sigmoid_prime = 18'b000000000001101001;
		14'b11000001011101:	sigmoid_prime = 18'b000000000001101001;
		14'b11000001011110:	sigmoid_prime = 18'b000000000001101001;
		14'b11000001011111:	sigmoid_prime = 18'b000000000001101001;
		14'b11000001100000:	sigmoid_prime = 18'b000000000001101001;
		14'b11000001100001:	sigmoid_prime = 18'b000000000001101010;
		14'b11000001100010:	sigmoid_prime = 18'b000000000001101010;
		14'b11000001100011:	sigmoid_prime = 18'b000000000001101010;
		14'b11000001100100:	sigmoid_prime = 18'b000000000001101010;
		14'b11000001100101:	sigmoid_prime = 18'b000000000001101011;
		14'b11000001100110:	sigmoid_prime = 18'b000000000001101011;
		14'b11000001100111:	sigmoid_prime = 18'b000000000001101011;
		14'b11000001101000:	sigmoid_prime = 18'b000000000001101011;
		14'b11000001101001:	sigmoid_prime = 18'b000000000001101011;
		14'b11000001101010:	sigmoid_prime = 18'b000000000001101100;
		14'b11000001101011:	sigmoid_prime = 18'b000000000001101100;
		14'b11000001101100:	sigmoid_prime = 18'b000000000001101100;
		14'b11000001101101:	sigmoid_prime = 18'b000000000001101100;
		14'b11000001101110:	sigmoid_prime = 18'b000000000001101100;
		14'b11000001101111:	sigmoid_prime = 18'b000000000001101101;
		14'b11000001110000:	sigmoid_prime = 18'b000000000001101101;
		14'b11000001110001:	sigmoid_prime = 18'b000000000001101101;
		14'b11000001110010:	sigmoid_prime = 18'b000000000001101101;
		14'b11000001110011:	sigmoid_prime = 18'b000000000001101101;
		14'b11000001110100:	sigmoid_prime = 18'b000000000001101110;
		14'b11000001110101:	sigmoid_prime = 18'b000000000001101110;
		14'b11000001110110:	sigmoid_prime = 18'b000000000001101110;
		14'b11000001110111:	sigmoid_prime = 18'b000000000001101110;
		14'b11000001111000:	sigmoid_prime = 18'b000000000001101111;
		14'b11000001111001:	sigmoid_prime = 18'b000000000001101111;
		14'b11000001111010:	sigmoid_prime = 18'b000000000001101111;
		14'b11000001111011:	sigmoid_prime = 18'b000000000001101111;
		14'b11000001111100:	sigmoid_prime = 18'b000000000001101111;
		14'b11000001111101:	sigmoid_prime = 18'b000000000001110000;
		14'b11000001111110:	sigmoid_prime = 18'b000000000001110000;
		14'b11000001111111:	sigmoid_prime = 18'b000000000001110000;
		14'b11000010000000:	sigmoid_prime = 18'b000000000001110000;
		14'b11000010000001:	sigmoid_prime = 18'b000000000001110001;
		14'b11000010000010:	sigmoid_prime = 18'b000000000001110001;
		14'b11000010000011:	sigmoid_prime = 18'b000000000001110001;
		14'b11000010000100:	sigmoid_prime = 18'b000000000001110001;
		14'b11000010000101:	sigmoid_prime = 18'b000000000001110001;
		14'b11000010000110:	sigmoid_prime = 18'b000000000001110010;
		14'b11000010000111:	sigmoid_prime = 18'b000000000001110010;
		14'b11000010001000:	sigmoid_prime = 18'b000000000001110010;
		14'b11000010001001:	sigmoid_prime = 18'b000000000001110010;
		14'b11000010001010:	sigmoid_prime = 18'b000000000001110011;
		14'b11000010001011:	sigmoid_prime = 18'b000000000001110011;
		14'b11000010001100:	sigmoid_prime = 18'b000000000001110011;
		14'b11000010001101:	sigmoid_prime = 18'b000000000001110011;
		14'b11000010001110:	sigmoid_prime = 18'b000000000001110011;
		14'b11000010001111:	sigmoid_prime = 18'b000000000001110100;
		14'b11000010010000:	sigmoid_prime = 18'b000000000001110100;
		14'b11000010010001:	sigmoid_prime = 18'b000000000001110100;
		14'b11000010010010:	sigmoid_prime = 18'b000000000001110100;
		14'b11000010010011:	sigmoid_prime = 18'b000000000001110101;
		14'b11000010010100:	sigmoid_prime = 18'b000000000001110101;
		14'b11000010010101:	sigmoid_prime = 18'b000000000001110101;
		14'b11000010010110:	sigmoid_prime = 18'b000000000001110101;
		14'b11000010010111:	sigmoid_prime = 18'b000000000001110101;
		14'b11000010011000:	sigmoid_prime = 18'b000000000001110110;
		14'b11000010011001:	sigmoid_prime = 18'b000000000001110110;
		14'b11000010011010:	sigmoid_prime = 18'b000000000001110110;
		14'b11000010011011:	sigmoid_prime = 18'b000000000001110110;
		14'b11000010011100:	sigmoid_prime = 18'b000000000001110111;
		14'b11000010011101:	sigmoid_prime = 18'b000000000001110111;
		14'b11000010011110:	sigmoid_prime = 18'b000000000001110111;
		14'b11000010011111:	sigmoid_prime = 18'b000000000001110111;
		14'b11000010100000:	sigmoid_prime = 18'b000000000001111000;
		14'b11000010100001:	sigmoid_prime = 18'b000000000001111000;
		14'b11000010100010:	sigmoid_prime = 18'b000000000001111000;
		14'b11000010100011:	sigmoid_prime = 18'b000000000001111000;
		14'b11000010100100:	sigmoid_prime = 18'b000000000001111001;
		14'b11000010100101:	sigmoid_prime = 18'b000000000001111001;
		14'b11000010100110:	sigmoid_prime = 18'b000000000001111001;
		14'b11000010100111:	sigmoid_prime = 18'b000000000001111001;
		14'b11000010101000:	sigmoid_prime = 18'b000000000001111001;
		14'b11000010101001:	sigmoid_prime = 18'b000000000001111010;
		14'b11000010101010:	sigmoid_prime = 18'b000000000001111010;
		14'b11000010101011:	sigmoid_prime = 18'b000000000001111010;
		14'b11000010101100:	sigmoid_prime = 18'b000000000001111010;
		14'b11000010101101:	sigmoid_prime = 18'b000000000001111011;
		14'b11000010101110:	sigmoid_prime = 18'b000000000001111011;
		14'b11000010101111:	sigmoid_prime = 18'b000000000001111011;
		14'b11000010110000:	sigmoid_prime = 18'b000000000001111011;
		14'b11000010110001:	sigmoid_prime = 18'b000000000001111100;
		14'b11000010110010:	sigmoid_prime = 18'b000000000001111100;
		14'b11000010110011:	sigmoid_prime = 18'b000000000001111100;
		14'b11000010110100:	sigmoid_prime = 18'b000000000001111100;
		14'b11000010110101:	sigmoid_prime = 18'b000000000001111101;
		14'b11000010110110:	sigmoid_prime = 18'b000000000001111101;
		14'b11000010110111:	sigmoid_prime = 18'b000000000001111101;
		14'b11000010111000:	sigmoid_prime = 18'b000000000001111101;
		14'b11000010111001:	sigmoid_prime = 18'b000000000001111110;
		14'b11000010111010:	sigmoid_prime = 18'b000000000001111110;
		14'b11000010111011:	sigmoid_prime = 18'b000000000001111110;
		14'b11000010111100:	sigmoid_prime = 18'b000000000001111110;
		14'b11000010111101:	sigmoid_prime = 18'b000000000001111111;
		14'b11000010111110:	sigmoid_prime = 18'b000000000001111111;
		14'b11000010111111:	sigmoid_prime = 18'b000000000001111111;
		14'b11000011000000:	sigmoid_prime = 18'b000000000001111111;
		14'b11000011000001:	sigmoid_prime = 18'b000000000010000000;
		14'b11000011000010:	sigmoid_prime = 18'b000000000010000000;
		14'b11000011000011:	sigmoid_prime = 18'b000000000010000000;
		14'b11000011000100:	sigmoid_prime = 18'b000000000010000000;
		14'b11000011000101:	sigmoid_prime = 18'b000000000010000001;
		14'b11000011000110:	sigmoid_prime = 18'b000000000010000001;
		14'b11000011000111:	sigmoid_prime = 18'b000000000010000001;
		14'b11000011001000:	sigmoid_prime = 18'b000000000010000001;
		14'b11000011001001:	sigmoid_prime = 18'b000000000010000010;
		14'b11000011001010:	sigmoid_prime = 18'b000000000010000010;
		14'b11000011001011:	sigmoid_prime = 18'b000000000010000010;
		14'b11000011001100:	sigmoid_prime = 18'b000000000010000010;
		14'b11000011001101:	sigmoid_prime = 18'b000000000010000011;
		14'b11000011001110:	sigmoid_prime = 18'b000000000010000011;
		14'b11000011001111:	sigmoid_prime = 18'b000000000010000011;
		14'b11000011010000:	sigmoid_prime = 18'b000000000010000011;
		14'b11000011010001:	sigmoid_prime = 18'b000000000010000100;
		14'b11000011010010:	sigmoid_prime = 18'b000000000010000100;
		14'b11000011010011:	sigmoid_prime = 18'b000000000010000100;
		14'b11000011010100:	sigmoid_prime = 18'b000000000010000100;
		14'b11000011010101:	sigmoid_prime = 18'b000000000010000101;
		14'b11000011010110:	sigmoid_prime = 18'b000000000010000101;
		14'b11000011010111:	sigmoid_prime = 18'b000000000010000101;
		14'b11000011011000:	sigmoid_prime = 18'b000000000010000101;
		14'b11000011011001:	sigmoid_prime = 18'b000000000010000110;
		14'b11000011011010:	sigmoid_prime = 18'b000000000010000110;
		14'b11000011011011:	sigmoid_prime = 18'b000000000010000110;
		14'b11000011011100:	sigmoid_prime = 18'b000000000010000111;
		14'b11000011011101:	sigmoid_prime = 18'b000000000010000111;
		14'b11000011011110:	sigmoid_prime = 18'b000000000010000111;
		14'b11000011011111:	sigmoid_prime = 18'b000000000010000111;
		14'b11000011100000:	sigmoid_prime = 18'b000000000010001000;
		14'b11000011100001:	sigmoid_prime = 18'b000000000010001000;
		14'b11000011100010:	sigmoid_prime = 18'b000000000010001000;
		14'b11000011100011:	sigmoid_prime = 18'b000000000010001000;
		14'b11000011100100:	sigmoid_prime = 18'b000000000010001001;
		14'b11000011100101:	sigmoid_prime = 18'b000000000010001001;
		14'b11000011100110:	sigmoid_prime = 18'b000000000010001001;
		14'b11000011100111:	sigmoid_prime = 18'b000000000010001001;
		14'b11000011101000:	sigmoid_prime = 18'b000000000010001010;
		14'b11000011101001:	sigmoid_prime = 18'b000000000010001010;
		14'b11000011101010:	sigmoid_prime = 18'b000000000010001010;
		14'b11000011101011:	sigmoid_prime = 18'b000000000010001011;
		14'b11000011101100:	sigmoid_prime = 18'b000000000010001011;
		14'b11000011101101:	sigmoid_prime = 18'b000000000010001011;
		14'b11000011101110:	sigmoid_prime = 18'b000000000010001011;
		14'b11000011101111:	sigmoid_prime = 18'b000000000010001100;
		14'b11000011110000:	sigmoid_prime = 18'b000000000010001100;
		14'b11000011110001:	sigmoid_prime = 18'b000000000010001100;
		14'b11000011110010:	sigmoid_prime = 18'b000000000010001100;
		14'b11000011110011:	sigmoid_prime = 18'b000000000010001101;
		14'b11000011110100:	sigmoid_prime = 18'b000000000010001101;
		14'b11000011110101:	sigmoid_prime = 18'b000000000010001101;
		14'b11000011110110:	sigmoid_prime = 18'b000000000010001110;
		14'b11000011110111:	sigmoid_prime = 18'b000000000010001110;
		14'b11000011111000:	sigmoid_prime = 18'b000000000010001110;
		14'b11000011111001:	sigmoid_prime = 18'b000000000010001110;
		14'b11000011111010:	sigmoid_prime = 18'b000000000010001111;
		14'b11000011111011:	sigmoid_prime = 18'b000000000010001111;
		14'b11000011111100:	sigmoid_prime = 18'b000000000010001111;
		14'b11000011111101:	sigmoid_prime = 18'b000000000010001111;
		14'b11000011111110:	sigmoid_prime = 18'b000000000010010000;
		14'b11000011111111:	sigmoid_prime = 18'b000000000010010000;
		14'b11000100000000:	sigmoid_prime = 18'b000000000010010000;
		14'b11000100000001:	sigmoid_prime = 18'b000000000010010001;
		14'b11000100000010:	sigmoid_prime = 18'b000000000010010001;
		14'b11000100000011:	sigmoid_prime = 18'b000000000010010001;
		14'b11000100000100:	sigmoid_prime = 18'b000000000010010001;
		14'b11000100000101:	sigmoid_prime = 18'b000000000010010010;
		14'b11000100000110:	sigmoid_prime = 18'b000000000010010010;
		14'b11000100000111:	sigmoid_prime = 18'b000000000010010010;
		14'b11000100001000:	sigmoid_prime = 18'b000000000010010011;
		14'b11000100001001:	sigmoid_prime = 18'b000000000010010011;
		14'b11000100001010:	sigmoid_prime = 18'b000000000010010011;
		14'b11000100001011:	sigmoid_prime = 18'b000000000010010011;
		14'b11000100001100:	sigmoid_prime = 18'b000000000010010100;
		14'b11000100001101:	sigmoid_prime = 18'b000000000010010100;
		14'b11000100001110:	sigmoid_prime = 18'b000000000010010100;
		14'b11000100001111:	sigmoid_prime = 18'b000000000010010101;
		14'b11000100010000:	sigmoid_prime = 18'b000000000010010101;
		14'b11000100010001:	sigmoid_prime = 18'b000000000010010101;
		14'b11000100010010:	sigmoid_prime = 18'b000000000010010110;
		14'b11000100010011:	sigmoid_prime = 18'b000000000010010110;
		14'b11000100010100:	sigmoid_prime = 18'b000000000010010110;
		14'b11000100010101:	sigmoid_prime = 18'b000000000010010110;
		14'b11000100010110:	sigmoid_prime = 18'b000000000010010111;
		14'b11000100010111:	sigmoid_prime = 18'b000000000010010111;
		14'b11000100011000:	sigmoid_prime = 18'b000000000010010111;
		14'b11000100011001:	sigmoid_prime = 18'b000000000010011000;
		14'b11000100011010:	sigmoid_prime = 18'b000000000010011000;
		14'b11000100011011:	sigmoid_prime = 18'b000000000010011000;
		14'b11000100011100:	sigmoid_prime = 18'b000000000010011000;
		14'b11000100011101:	sigmoid_prime = 18'b000000000010011001;
		14'b11000100011110:	sigmoid_prime = 18'b000000000010011001;
		14'b11000100011111:	sigmoid_prime = 18'b000000000010011001;
		14'b11000100100000:	sigmoid_prime = 18'b000000000010011010;
		14'b11000100100001:	sigmoid_prime = 18'b000000000010011010;
		14'b11000100100010:	sigmoid_prime = 18'b000000000010011010;
		14'b11000100100011:	sigmoid_prime = 18'b000000000010011011;
		14'b11000100100100:	sigmoid_prime = 18'b000000000010011011;
		14'b11000100100101:	sigmoid_prime = 18'b000000000010011011;
		14'b11000100100110:	sigmoid_prime = 18'b000000000010011011;
		14'b11000100100111:	sigmoid_prime = 18'b000000000010011100;
		14'b11000100101000:	sigmoid_prime = 18'b000000000010011100;
		14'b11000100101001:	sigmoid_prime = 18'b000000000010011100;
		14'b11000100101010:	sigmoid_prime = 18'b000000000010011101;
		14'b11000100101011:	sigmoid_prime = 18'b000000000010011101;
		14'b11000100101100:	sigmoid_prime = 18'b000000000010011101;
		14'b11000100101101:	sigmoid_prime = 18'b000000000010011110;
		14'b11000100101110:	sigmoid_prime = 18'b000000000010011110;
		14'b11000100101111:	sigmoid_prime = 18'b000000000010011110;
		14'b11000100110000:	sigmoid_prime = 18'b000000000010011111;
		14'b11000100110001:	sigmoid_prime = 18'b000000000010011111;
		14'b11000100110010:	sigmoid_prime = 18'b000000000010011111;
		14'b11000100110011:	sigmoid_prime = 18'b000000000010011111;
		14'b11000100110100:	sigmoid_prime = 18'b000000000010100000;
		14'b11000100110101:	sigmoid_prime = 18'b000000000010100000;
		14'b11000100110110:	sigmoid_prime = 18'b000000000010100000;
		14'b11000100110111:	sigmoid_prime = 18'b000000000010100001;
		14'b11000100111000:	sigmoid_prime = 18'b000000000010100001;
		14'b11000100111001:	sigmoid_prime = 18'b000000000010100001;
		14'b11000100111010:	sigmoid_prime = 18'b000000000010100010;
		14'b11000100111011:	sigmoid_prime = 18'b000000000010100010;
		14'b11000100111100:	sigmoid_prime = 18'b000000000010100010;
		14'b11000100111101:	sigmoid_prime = 18'b000000000010100011;
		14'b11000100111110:	sigmoid_prime = 18'b000000000010100011;
		14'b11000100111111:	sigmoid_prime = 18'b000000000010100011;
		14'b11000101000000:	sigmoid_prime = 18'b000000000010100100;
		14'b11000101000001:	sigmoid_prime = 18'b000000000010100100;
		14'b11000101000010:	sigmoid_prime = 18'b000000000010100100;
		14'b11000101000011:	sigmoid_prime = 18'b000000000010100101;
		14'b11000101000100:	sigmoid_prime = 18'b000000000010100101;
		14'b11000101000101:	sigmoid_prime = 18'b000000000010100101;
		14'b11000101000110:	sigmoid_prime = 18'b000000000010100110;
		14'b11000101000111:	sigmoid_prime = 18'b000000000010100110;
		14'b11000101001000:	sigmoid_prime = 18'b000000000010100110;
		14'b11000101001001:	sigmoid_prime = 18'b000000000010100110;
		14'b11000101001010:	sigmoid_prime = 18'b000000000010100111;
		14'b11000101001011:	sigmoid_prime = 18'b000000000010100111;
		14'b11000101001100:	sigmoid_prime = 18'b000000000010100111;
		14'b11000101001101:	sigmoid_prime = 18'b000000000010101000;
		14'b11000101001110:	sigmoid_prime = 18'b000000000010101000;
		14'b11000101001111:	sigmoid_prime = 18'b000000000010101000;
		14'b11000101010000:	sigmoid_prime = 18'b000000000010101001;
		14'b11000101010001:	sigmoid_prime = 18'b000000000010101001;
		14'b11000101010010:	sigmoid_prime = 18'b000000000010101001;
		14'b11000101010011:	sigmoid_prime = 18'b000000000010101010;
		14'b11000101010100:	sigmoid_prime = 18'b000000000010101010;
		14'b11000101010101:	sigmoid_prime = 18'b000000000010101010;
		14'b11000101010110:	sigmoid_prime = 18'b000000000010101011;
		14'b11000101010111:	sigmoid_prime = 18'b000000000010101011;
		14'b11000101011000:	sigmoid_prime = 18'b000000000010101011;
		14'b11000101011001:	sigmoid_prime = 18'b000000000010101100;
		14'b11000101011010:	sigmoid_prime = 18'b000000000010101100;
		14'b11000101011011:	sigmoid_prime = 18'b000000000010101100;
		14'b11000101011100:	sigmoid_prime = 18'b000000000010101101;
		14'b11000101011101:	sigmoid_prime = 18'b000000000010101101;
		14'b11000101011110:	sigmoid_prime = 18'b000000000010101101;
		14'b11000101011111:	sigmoid_prime = 18'b000000000010101110;
		14'b11000101100000:	sigmoid_prime = 18'b000000000010101110;
		14'b11000101100001:	sigmoid_prime = 18'b000000000010101110;
		14'b11000101100010:	sigmoid_prime = 18'b000000000010101111;
		14'b11000101100011:	sigmoid_prime = 18'b000000000010101111;
		14'b11000101100100:	sigmoid_prime = 18'b000000000010110000;
		14'b11000101100101:	sigmoid_prime = 18'b000000000010110000;
		14'b11000101100110:	sigmoid_prime = 18'b000000000010110000;
		14'b11000101100111:	sigmoid_prime = 18'b000000000010110001;
		14'b11000101101000:	sigmoid_prime = 18'b000000000010110001;
		14'b11000101101001:	sigmoid_prime = 18'b000000000010110001;
		14'b11000101101010:	sigmoid_prime = 18'b000000000010110010;
		14'b11000101101011:	sigmoid_prime = 18'b000000000010110010;
		14'b11000101101100:	sigmoid_prime = 18'b000000000010110010;
		14'b11000101101101:	sigmoid_prime = 18'b000000000010110011;
		14'b11000101101110:	sigmoid_prime = 18'b000000000010110011;
		14'b11000101101111:	sigmoid_prime = 18'b000000000010110011;
		14'b11000101110000:	sigmoid_prime = 18'b000000000010110100;
		14'b11000101110001:	sigmoid_prime = 18'b000000000010110100;
		14'b11000101110010:	sigmoid_prime = 18'b000000000010110100;
		14'b11000101110011:	sigmoid_prime = 18'b000000000010110101;
		14'b11000101110100:	sigmoid_prime = 18'b000000000010110101;
		14'b11000101110101:	sigmoid_prime = 18'b000000000010110101;
		14'b11000101110110:	sigmoid_prime = 18'b000000000010110110;
		14'b11000101110111:	sigmoid_prime = 18'b000000000010110110;
		14'b11000101111000:	sigmoid_prime = 18'b000000000010110111;
		14'b11000101111001:	sigmoid_prime = 18'b000000000010110111;
		14'b11000101111010:	sigmoid_prime = 18'b000000000010110111;
		14'b11000101111011:	sigmoid_prime = 18'b000000000010111000;
		14'b11000101111100:	sigmoid_prime = 18'b000000000010111000;
		14'b11000101111101:	sigmoid_prime = 18'b000000000010111000;
		14'b11000101111110:	sigmoid_prime = 18'b000000000010111001;
		14'b11000101111111:	sigmoid_prime = 18'b000000000010111001;
		14'b11000110000000:	sigmoid_prime = 18'b000000000010111001;
		14'b11000110000001:	sigmoid_prime = 18'b000000000010111010;
		14'b11000110000010:	sigmoid_prime = 18'b000000000010111010;
		14'b11000110000011:	sigmoid_prime = 18'b000000000010111010;
		14'b11000110000100:	sigmoid_prime = 18'b000000000010111011;
		14'b11000110000101:	sigmoid_prime = 18'b000000000010111011;
		14'b11000110000110:	sigmoid_prime = 18'b000000000010111100;
		14'b11000110000111:	sigmoid_prime = 18'b000000000010111100;
		14'b11000110001000:	sigmoid_prime = 18'b000000000010111100;
		14'b11000110001001:	sigmoid_prime = 18'b000000000010111101;
		14'b11000110001010:	sigmoid_prime = 18'b000000000010111101;
		14'b11000110001011:	sigmoid_prime = 18'b000000000010111101;
		14'b11000110001100:	sigmoid_prime = 18'b000000000010111110;
		14'b11000110001101:	sigmoid_prime = 18'b000000000010111110;
		14'b11000110001110:	sigmoid_prime = 18'b000000000010111111;
		14'b11000110001111:	sigmoid_prime = 18'b000000000010111111;
		14'b11000110010000:	sigmoid_prime = 18'b000000000010111111;
		14'b11000110010001:	sigmoid_prime = 18'b000000000011000000;
		14'b11000110010010:	sigmoid_prime = 18'b000000000011000000;
		14'b11000110010011:	sigmoid_prime = 18'b000000000011000000;
		14'b11000110010100:	sigmoid_prime = 18'b000000000011000001;
		14'b11000110010101:	sigmoid_prime = 18'b000000000011000001;
		14'b11000110010110:	sigmoid_prime = 18'b000000000011000010;
		14'b11000110010111:	sigmoid_prime = 18'b000000000011000010;
		14'b11000110011000:	sigmoid_prime = 18'b000000000011000010;
		14'b11000110011001:	sigmoid_prime = 18'b000000000011000011;
		14'b11000110011010:	sigmoid_prime = 18'b000000000011000011;
		14'b11000110011011:	sigmoid_prime = 18'b000000000011000011;
		14'b11000110011100:	sigmoid_prime = 18'b000000000011000100;
		14'b11000110011101:	sigmoid_prime = 18'b000000000011000100;
		14'b11000110011110:	sigmoid_prime = 18'b000000000011000101;
		14'b11000110011111:	sigmoid_prime = 18'b000000000011000101;
		14'b11000110100000:	sigmoid_prime = 18'b000000000011000101;
		14'b11000110100001:	sigmoid_prime = 18'b000000000011000110;
		14'b11000110100010:	sigmoid_prime = 18'b000000000011000110;
		14'b11000110100011:	sigmoid_prime = 18'b000000000011000111;
		14'b11000110100100:	sigmoid_prime = 18'b000000000011000111;
		14'b11000110100101:	sigmoid_prime = 18'b000000000011000111;
		14'b11000110100110:	sigmoid_prime = 18'b000000000011001000;
		14'b11000110100111:	sigmoid_prime = 18'b000000000011001000;
		14'b11000110101000:	sigmoid_prime = 18'b000000000011001000;
		14'b11000110101001:	sigmoid_prime = 18'b000000000011001001;
		14'b11000110101010:	sigmoid_prime = 18'b000000000011001001;
		14'b11000110101011:	sigmoid_prime = 18'b000000000011001010;
		14'b11000110101100:	sigmoid_prime = 18'b000000000011001010;
		14'b11000110101101:	sigmoid_prime = 18'b000000000011001010;
		14'b11000110101110:	sigmoid_prime = 18'b000000000011001011;
		14'b11000110101111:	sigmoid_prime = 18'b000000000011001011;
		14'b11000110110000:	sigmoid_prime = 18'b000000000011001100;
		14'b11000110110001:	sigmoid_prime = 18'b000000000011001100;
		14'b11000110110010:	sigmoid_prime = 18'b000000000011001100;
		14'b11000110110011:	sigmoid_prime = 18'b000000000011001101;
		14'b11000110110100:	sigmoid_prime = 18'b000000000011001101;
		14'b11000110110101:	sigmoid_prime = 18'b000000000011001110;
		14'b11000110110110:	sigmoid_prime = 18'b000000000011001110;
		14'b11000110110111:	sigmoid_prime = 18'b000000000011001110;
		14'b11000110111000:	sigmoid_prime = 18'b000000000011001111;
		14'b11000110111001:	sigmoid_prime = 18'b000000000011001111;
		14'b11000110111010:	sigmoid_prime = 18'b000000000011010000;
		14'b11000110111011:	sigmoid_prime = 18'b000000000011010000;
		14'b11000110111100:	sigmoid_prime = 18'b000000000011010000;
		14'b11000110111101:	sigmoid_prime = 18'b000000000011010001;
		14'b11000110111110:	sigmoid_prime = 18'b000000000011010001;
		14'b11000110111111:	sigmoid_prime = 18'b000000000011010010;
		14'b11000111000000:	sigmoid_prime = 18'b000000000011010010;
		14'b11000111000001:	sigmoid_prime = 18'b000000000011010011;
		14'b11000111000010:	sigmoid_prime = 18'b000000000011010011;
		14'b11000111000011:	sigmoid_prime = 18'b000000000011010011;
		14'b11000111000100:	sigmoid_prime = 18'b000000000011010100;
		14'b11000111000101:	sigmoid_prime = 18'b000000000011010100;
		14'b11000111000110:	sigmoid_prime = 18'b000000000011010101;
		14'b11000111000111:	sigmoid_prime = 18'b000000000011010101;
		14'b11000111001000:	sigmoid_prime = 18'b000000000011010101;
		14'b11000111001001:	sigmoid_prime = 18'b000000000011010110;
		14'b11000111001010:	sigmoid_prime = 18'b000000000011010110;
		14'b11000111001011:	sigmoid_prime = 18'b000000000011010111;
		14'b11000111001100:	sigmoid_prime = 18'b000000000011010111;
		14'b11000111001101:	sigmoid_prime = 18'b000000000011011000;
		14'b11000111001110:	sigmoid_prime = 18'b000000000011011000;
		14'b11000111001111:	sigmoid_prime = 18'b000000000011011000;
		14'b11000111010000:	sigmoid_prime = 18'b000000000011011001;
		14'b11000111010001:	sigmoid_prime = 18'b000000000011011001;
		14'b11000111010010:	sigmoid_prime = 18'b000000000011011010;
		14'b11000111010011:	sigmoid_prime = 18'b000000000011011010;
		14'b11000111010100:	sigmoid_prime = 18'b000000000011011010;
		14'b11000111010101:	sigmoid_prime = 18'b000000000011011011;
		14'b11000111010110:	sigmoid_prime = 18'b000000000011011011;
		14'b11000111010111:	sigmoid_prime = 18'b000000000011011100;
		14'b11000111011000:	sigmoid_prime = 18'b000000000011011100;
		14'b11000111011001:	sigmoid_prime = 18'b000000000011011101;
		14'b11000111011010:	sigmoid_prime = 18'b000000000011011101;
		14'b11000111011011:	sigmoid_prime = 18'b000000000011011110;
		14'b11000111011100:	sigmoid_prime = 18'b000000000011011110;
		14'b11000111011101:	sigmoid_prime = 18'b000000000011011110;
		14'b11000111011110:	sigmoid_prime = 18'b000000000011011111;
		14'b11000111011111:	sigmoid_prime = 18'b000000000011011111;
		14'b11000111100000:	sigmoid_prime = 18'b000000000011100000;
		14'b11000111100001:	sigmoid_prime = 18'b000000000011100000;
		14'b11000111100010:	sigmoid_prime = 18'b000000000011100001;
		14'b11000111100011:	sigmoid_prime = 18'b000000000011100001;
		14'b11000111100100:	sigmoid_prime = 18'b000000000011100001;
		14'b11000111100101:	sigmoid_prime = 18'b000000000011100010;
		14'b11000111100110:	sigmoid_prime = 18'b000000000011100010;
		14'b11000111100111:	sigmoid_prime = 18'b000000000011100011;
		14'b11000111101000:	sigmoid_prime = 18'b000000000011100011;
		14'b11000111101001:	sigmoid_prime = 18'b000000000011100100;
		14'b11000111101010:	sigmoid_prime = 18'b000000000011100100;
		14'b11000111101011:	sigmoid_prime = 18'b000000000011100101;
		14'b11000111101100:	sigmoid_prime = 18'b000000000011100101;
		14'b11000111101101:	sigmoid_prime = 18'b000000000011100101;
		14'b11000111101110:	sigmoid_prime = 18'b000000000011100110;
		14'b11000111101111:	sigmoid_prime = 18'b000000000011100110;
		14'b11000111110000:	sigmoid_prime = 18'b000000000011100111;
		14'b11000111110001:	sigmoid_prime = 18'b000000000011100111;
		14'b11000111110010:	sigmoid_prime = 18'b000000000011101000;
		14'b11000111110011:	sigmoid_prime = 18'b000000000011101000;
		14'b11000111110100:	sigmoid_prime = 18'b000000000011101001;
		14'b11000111110101:	sigmoid_prime = 18'b000000000011101001;
		14'b11000111110110:	sigmoid_prime = 18'b000000000011101010;
		14'b11000111110111:	sigmoid_prime = 18'b000000000011101010;
		14'b11000111111000:	sigmoid_prime = 18'b000000000011101010;
		14'b11000111111001:	sigmoid_prime = 18'b000000000011101011;
		14'b11000111111010:	sigmoid_prime = 18'b000000000011101011;
		14'b11000111111011:	sigmoid_prime = 18'b000000000011101100;
		14'b11000111111100:	sigmoid_prime = 18'b000000000011101100;
		14'b11000111111101:	sigmoid_prime = 18'b000000000011101101;
		14'b11000111111110:	sigmoid_prime = 18'b000000000011101101;
		14'b11000111111111:	sigmoid_prime = 18'b000000000011101110;
		14'b11001000000000:	sigmoid_prime = 18'b000000000011101110;
		14'b11001000000001:	sigmoid_prime = 18'b000000000011101111;
		14'b11001000000010:	sigmoid_prime = 18'b000000000011101111;
		14'b11001000000011:	sigmoid_prime = 18'b000000000011110000;
		14'b11001000000100:	sigmoid_prime = 18'b000000000011110000;
		14'b11001000000101:	sigmoid_prime = 18'b000000000011110000;
		14'b11001000000110:	sigmoid_prime = 18'b000000000011110001;
		14'b11001000000111:	sigmoid_prime = 18'b000000000011110001;
		14'b11001000001000:	sigmoid_prime = 18'b000000000011110010;
		14'b11001000001001:	sigmoid_prime = 18'b000000000011110010;
		14'b11001000001010:	sigmoid_prime = 18'b000000000011110011;
		14'b11001000001011:	sigmoid_prime = 18'b000000000011110011;
		14'b11001000001100:	sigmoid_prime = 18'b000000000011110100;
		14'b11001000001101:	sigmoid_prime = 18'b000000000011110100;
		14'b11001000001110:	sigmoid_prime = 18'b000000000011110101;
		14'b11001000001111:	sigmoid_prime = 18'b000000000011110101;
		14'b11001000010000:	sigmoid_prime = 18'b000000000011110110;
		14'b11001000010001:	sigmoid_prime = 18'b000000000011110110;
		14'b11001000010010:	sigmoid_prime = 18'b000000000011110111;
		14'b11001000010011:	sigmoid_prime = 18'b000000000011110111;
		14'b11001000010100:	sigmoid_prime = 18'b000000000011111000;
		14'b11001000010101:	sigmoid_prime = 18'b000000000011111000;
		14'b11001000010110:	sigmoid_prime = 18'b000000000011111001;
		14'b11001000010111:	sigmoid_prime = 18'b000000000011111001;
		14'b11001000011000:	sigmoid_prime = 18'b000000000011111010;
		14'b11001000011001:	sigmoid_prime = 18'b000000000011111010;
		14'b11001000011010:	sigmoid_prime = 18'b000000000011111011;
		14'b11001000011011:	sigmoid_prime = 18'b000000000011111011;
		14'b11001000011100:	sigmoid_prime = 18'b000000000011111011;
		14'b11001000011101:	sigmoid_prime = 18'b000000000011111100;
		14'b11001000011110:	sigmoid_prime = 18'b000000000011111100;
		14'b11001000011111:	sigmoid_prime = 18'b000000000011111101;
		14'b11001000100000:	sigmoid_prime = 18'b000000000011111101;
		14'b11001000100001:	sigmoid_prime = 18'b000000000011111110;
		14'b11001000100010:	sigmoid_prime = 18'b000000000011111110;
		14'b11001000100011:	sigmoid_prime = 18'b000000000011111111;
		14'b11001000100100:	sigmoid_prime = 18'b000000000011111111;
		14'b11001000100101:	sigmoid_prime = 18'b000000000100000000;
		14'b11001000100110:	sigmoid_prime = 18'b000000000100000000;
		14'b11001000100111:	sigmoid_prime = 18'b000000000100000001;
		14'b11001000101000:	sigmoid_prime = 18'b000000000100000001;
		14'b11001000101001:	sigmoid_prime = 18'b000000000100000010;
		14'b11001000101010:	sigmoid_prime = 18'b000000000100000010;
		14'b11001000101011:	sigmoid_prime = 18'b000000000100000011;
		14'b11001000101100:	sigmoid_prime = 18'b000000000100000011;
		14'b11001000101101:	sigmoid_prime = 18'b000000000100000100;
		14'b11001000101110:	sigmoid_prime = 18'b000000000100000100;
		14'b11001000101111:	sigmoid_prime = 18'b000000000100000101;
		14'b11001000110000:	sigmoid_prime = 18'b000000000100000110;
		14'b11001000110001:	sigmoid_prime = 18'b000000000100000110;
		14'b11001000110010:	sigmoid_prime = 18'b000000000100000111;
		14'b11001000110011:	sigmoid_prime = 18'b000000000100000111;
		14'b11001000110100:	sigmoid_prime = 18'b000000000100001000;
		14'b11001000110101:	sigmoid_prime = 18'b000000000100001000;
		14'b11001000110110:	sigmoid_prime = 18'b000000000100001001;
		14'b11001000110111:	sigmoid_prime = 18'b000000000100001001;
		14'b11001000111000:	sigmoid_prime = 18'b000000000100001010;
		14'b11001000111001:	sigmoid_prime = 18'b000000000100001010;
		14'b11001000111010:	sigmoid_prime = 18'b000000000100001011;
		14'b11001000111011:	sigmoid_prime = 18'b000000000100001011;
		14'b11001000111100:	sigmoid_prime = 18'b000000000100001100;
		14'b11001000111101:	sigmoid_prime = 18'b000000000100001100;
		14'b11001000111110:	sigmoid_prime = 18'b000000000100001101;
		14'b11001000111111:	sigmoid_prime = 18'b000000000100001101;
		14'b11001001000000:	sigmoid_prime = 18'b000000000100001110;
		14'b11001001000001:	sigmoid_prime = 18'b000000000100001110;
		14'b11001001000010:	sigmoid_prime = 18'b000000000100001111;
		14'b11001001000011:	sigmoid_prime = 18'b000000000100001111;
		14'b11001001000100:	sigmoid_prime = 18'b000000000100010000;
		14'b11001001000101:	sigmoid_prime = 18'b000000000100010000;
		14'b11001001000110:	sigmoid_prime = 18'b000000000100010001;
		14'b11001001000111:	sigmoid_prime = 18'b000000000100010010;
		14'b11001001001000:	sigmoid_prime = 18'b000000000100010010;
		14'b11001001001001:	sigmoid_prime = 18'b000000000100010011;
		14'b11001001001010:	sigmoid_prime = 18'b000000000100010011;
		14'b11001001001011:	sigmoid_prime = 18'b000000000100010100;
		14'b11001001001100:	sigmoid_prime = 18'b000000000100010100;
		14'b11001001001101:	sigmoid_prime = 18'b000000000100010101;
		14'b11001001001110:	sigmoid_prime = 18'b000000000100010101;
		14'b11001001001111:	sigmoid_prime = 18'b000000000100010110;
		14'b11001001010000:	sigmoid_prime = 18'b000000000100010110;
		14'b11001001010001:	sigmoid_prime = 18'b000000000100010111;
		14'b11001001010010:	sigmoid_prime = 18'b000000000100010111;
		14'b11001001010011:	sigmoid_prime = 18'b000000000100011000;
		14'b11001001010100:	sigmoid_prime = 18'b000000000100011001;
		14'b11001001010101:	sigmoid_prime = 18'b000000000100011001;
		14'b11001001010110:	sigmoid_prime = 18'b000000000100011010;
		14'b11001001010111:	sigmoid_prime = 18'b000000000100011010;
		14'b11001001011000:	sigmoid_prime = 18'b000000000100011011;
		14'b11001001011001:	sigmoid_prime = 18'b000000000100011011;
		14'b11001001011010:	sigmoid_prime = 18'b000000000100011100;
		14'b11001001011011:	sigmoid_prime = 18'b000000000100011100;
		14'b11001001011100:	sigmoid_prime = 18'b000000000100011101;
		14'b11001001011101:	sigmoid_prime = 18'b000000000100011110;
		14'b11001001011110:	sigmoid_prime = 18'b000000000100011110;
		14'b11001001011111:	sigmoid_prime = 18'b000000000100011111;
		14'b11001001100000:	sigmoid_prime = 18'b000000000100011111;
		14'b11001001100001:	sigmoid_prime = 18'b000000000100100000;
		14'b11001001100010:	sigmoid_prime = 18'b000000000100100000;
		14'b11001001100011:	sigmoid_prime = 18'b000000000100100001;
		14'b11001001100100:	sigmoid_prime = 18'b000000000100100001;
		14'b11001001100101:	sigmoid_prime = 18'b000000000100100010;
		14'b11001001100110:	sigmoid_prime = 18'b000000000100100011;
		14'b11001001100111:	sigmoid_prime = 18'b000000000100100011;
		14'b11001001101000:	sigmoid_prime = 18'b000000000100100100;
		14'b11001001101001:	sigmoid_prime = 18'b000000000100100100;
		14'b11001001101010:	sigmoid_prime = 18'b000000000100100101;
		14'b11001001101011:	sigmoid_prime = 18'b000000000100100101;
		14'b11001001101100:	sigmoid_prime = 18'b000000000100100110;
		14'b11001001101101:	sigmoid_prime = 18'b000000000100100111;
		14'b11001001101110:	sigmoid_prime = 18'b000000000100100111;
		14'b11001001101111:	sigmoid_prime = 18'b000000000100101000;
		14'b11001001110000:	sigmoid_prime = 18'b000000000100101000;
		14'b11001001110001:	sigmoid_prime = 18'b000000000100101001;
		14'b11001001110010:	sigmoid_prime = 18'b000000000100101001;
		14'b11001001110011:	sigmoid_prime = 18'b000000000100101010;
		14'b11001001110100:	sigmoid_prime = 18'b000000000100101011;
		14'b11001001110101:	sigmoid_prime = 18'b000000000100101011;
		14'b11001001110110:	sigmoid_prime = 18'b000000000100101100;
		14'b11001001110111:	sigmoid_prime = 18'b000000000100101100;
		14'b11001001111000:	sigmoid_prime = 18'b000000000100101101;
		14'b11001001111001:	sigmoid_prime = 18'b000000000100101110;
		14'b11001001111010:	sigmoid_prime = 18'b000000000100101110;
		14'b11001001111011:	sigmoid_prime = 18'b000000000100101111;
		14'b11001001111100:	sigmoid_prime = 18'b000000000100101111;
		14'b11001001111101:	sigmoid_prime = 18'b000000000100110000;
		14'b11001001111110:	sigmoid_prime = 18'b000000000100110001;
		14'b11001001111111:	sigmoid_prime = 18'b000000000100110001;
		14'b11001010000000:	sigmoid_prime = 18'b000000000100110010;
		14'b11001010000001:	sigmoid_prime = 18'b000000000100110010;
		14'b11001010000010:	sigmoid_prime = 18'b000000000100110011;
		14'b11001010000011:	sigmoid_prime = 18'b000000000100110100;
		14'b11001010000100:	sigmoid_prime = 18'b000000000100110100;
		14'b11001010000101:	sigmoid_prime = 18'b000000000100110101;
		14'b11001010000110:	sigmoid_prime = 18'b000000000100110101;
		14'b11001010000111:	sigmoid_prime = 18'b000000000100110110;
		14'b11001010001000:	sigmoid_prime = 18'b000000000100110111;
		14'b11001010001001:	sigmoid_prime = 18'b000000000100110111;
		14'b11001010001010:	sigmoid_prime = 18'b000000000100111000;
		14'b11001010001011:	sigmoid_prime = 18'b000000000100111000;
		14'b11001010001100:	sigmoid_prime = 18'b000000000100111001;
		14'b11001010001101:	sigmoid_prime = 18'b000000000100111010;
		14'b11001010001110:	sigmoid_prime = 18'b000000000100111010;
		14'b11001010001111:	sigmoid_prime = 18'b000000000100111011;
		14'b11001010010000:	sigmoid_prime = 18'b000000000100111011;
		14'b11001010010001:	sigmoid_prime = 18'b000000000100111100;
		14'b11001010010010:	sigmoid_prime = 18'b000000000100111101;
		14'b11001010010011:	sigmoid_prime = 18'b000000000100111101;
		14'b11001010010100:	sigmoid_prime = 18'b000000000100111110;
		14'b11001010010101:	sigmoid_prime = 18'b000000000100111111;
		14'b11001010010110:	sigmoid_prime = 18'b000000000100111111;
		14'b11001010010111:	sigmoid_prime = 18'b000000000101000000;
		14'b11001010011000:	sigmoid_prime = 18'b000000000101000000;
		14'b11001010011001:	sigmoid_prime = 18'b000000000101000001;
		14'b11001010011010:	sigmoid_prime = 18'b000000000101000010;
		14'b11001010011011:	sigmoid_prime = 18'b000000000101000010;
		14'b11001010011100:	sigmoid_prime = 18'b000000000101000011;
		14'b11001010011101:	sigmoid_prime = 18'b000000000101000100;
		14'b11001010011110:	sigmoid_prime = 18'b000000000101000100;
		14'b11001010011111:	sigmoid_prime = 18'b000000000101000101;
		14'b11001010100000:	sigmoid_prime = 18'b000000000101000101;
		14'b11001010100001:	sigmoid_prime = 18'b000000000101000110;
		14'b11001010100010:	sigmoid_prime = 18'b000000000101000111;
		14'b11001010100011:	sigmoid_prime = 18'b000000000101000111;
		14'b11001010100100:	sigmoid_prime = 18'b000000000101001000;
		14'b11001010100101:	sigmoid_prime = 18'b000000000101001001;
		14'b11001010100110:	sigmoid_prime = 18'b000000000101001001;
		14'b11001010100111:	sigmoid_prime = 18'b000000000101001010;
		14'b11001010101000:	sigmoid_prime = 18'b000000000101001011;
		14'b11001010101001:	sigmoid_prime = 18'b000000000101001011;
		14'b11001010101010:	sigmoid_prime = 18'b000000000101001100;
		14'b11001010101011:	sigmoid_prime = 18'b000000000101001100;
		14'b11001010101100:	sigmoid_prime = 18'b000000000101001101;
		14'b11001010101101:	sigmoid_prime = 18'b000000000101001110;
		14'b11001010101110:	sigmoid_prime = 18'b000000000101001110;
		14'b11001010101111:	sigmoid_prime = 18'b000000000101001111;
		14'b11001010110000:	sigmoid_prime = 18'b000000000101010000;
		14'b11001010110001:	sigmoid_prime = 18'b000000000101010000;
		14'b11001010110010:	sigmoid_prime = 18'b000000000101010001;
		14'b11001010110011:	sigmoid_prime = 18'b000000000101010010;
		14'b11001010110100:	sigmoid_prime = 18'b000000000101010010;
		14'b11001010110101:	sigmoid_prime = 18'b000000000101010011;
		14'b11001010110110:	sigmoid_prime = 18'b000000000101010100;
		14'b11001010110111:	sigmoid_prime = 18'b000000000101010100;
		14'b11001010111000:	sigmoid_prime = 18'b000000000101010101;
		14'b11001010111001:	sigmoid_prime = 18'b000000000101010110;
		14'b11001010111010:	sigmoid_prime = 18'b000000000101010110;
		14'b11001010111011:	sigmoid_prime = 18'b000000000101010111;
		14'b11001010111100:	sigmoid_prime = 18'b000000000101011000;
		14'b11001010111101:	sigmoid_prime = 18'b000000000101011000;
		14'b11001010111110:	sigmoid_prime = 18'b000000000101011001;
		14'b11001010111111:	sigmoid_prime = 18'b000000000101011010;
		14'b11001011000000:	sigmoid_prime = 18'b000000000101011010;
		14'b11001011000001:	sigmoid_prime = 18'b000000000101011011;
		14'b11001011000010:	sigmoid_prime = 18'b000000000101011100;
		14'b11001011000011:	sigmoid_prime = 18'b000000000101011100;
		14'b11001011000100:	sigmoid_prime = 18'b000000000101011101;
		14'b11001011000101:	sigmoid_prime = 18'b000000000101011110;
		14'b11001011000110:	sigmoid_prime = 18'b000000000101011110;
		14'b11001011000111:	sigmoid_prime = 18'b000000000101011111;
		14'b11001011001000:	sigmoid_prime = 18'b000000000101100000;
		14'b11001011001001:	sigmoid_prime = 18'b000000000101100001;
		14'b11001011001010:	sigmoid_prime = 18'b000000000101100001;
		14'b11001011001011:	sigmoid_prime = 18'b000000000101100010;
		14'b11001011001100:	sigmoid_prime = 18'b000000000101100011;
		14'b11001011001101:	sigmoid_prime = 18'b000000000101100011;
		14'b11001011001110:	sigmoid_prime = 18'b000000000101100100;
		14'b11001011001111:	sigmoid_prime = 18'b000000000101100101;
		14'b11001011010000:	sigmoid_prime = 18'b000000000101100101;
		14'b11001011010001:	sigmoid_prime = 18'b000000000101100110;
		14'b11001011010010:	sigmoid_prime = 18'b000000000101100111;
		14'b11001011010011:	sigmoid_prime = 18'b000000000101100111;
		14'b11001011010100:	sigmoid_prime = 18'b000000000101101000;
		14'b11001011010101:	sigmoid_prime = 18'b000000000101101001;
		14'b11001011010110:	sigmoid_prime = 18'b000000000101101010;
		14'b11001011010111:	sigmoid_prime = 18'b000000000101101010;
		14'b11001011011000:	sigmoid_prime = 18'b000000000101101011;
		14'b11001011011001:	sigmoid_prime = 18'b000000000101101100;
		14'b11001011011010:	sigmoid_prime = 18'b000000000101101100;
		14'b11001011011011:	sigmoid_prime = 18'b000000000101101101;
		14'b11001011011100:	sigmoid_prime = 18'b000000000101101110;
		14'b11001011011101:	sigmoid_prime = 18'b000000000101101111;
		14'b11001011011110:	sigmoid_prime = 18'b000000000101101111;
		14'b11001011011111:	sigmoid_prime = 18'b000000000101110000;
		14'b11001011100000:	sigmoid_prime = 18'b000000000101110001;
		14'b11001011100001:	sigmoid_prime = 18'b000000000101110001;
		14'b11001011100010:	sigmoid_prime = 18'b000000000101110010;
		14'b11001011100011:	sigmoid_prime = 18'b000000000101110011;
		14'b11001011100100:	sigmoid_prime = 18'b000000000101110100;
		14'b11001011100101:	sigmoid_prime = 18'b000000000101110100;
		14'b11001011100110:	sigmoid_prime = 18'b000000000101110101;
		14'b11001011100111:	sigmoid_prime = 18'b000000000101110110;
		14'b11001011101000:	sigmoid_prime = 18'b000000000101110110;
		14'b11001011101001:	sigmoid_prime = 18'b000000000101110111;
		14'b11001011101010:	sigmoid_prime = 18'b000000000101111000;
		14'b11001011101011:	sigmoid_prime = 18'b000000000101111001;
		14'b11001011101100:	sigmoid_prime = 18'b000000000101111001;
		14'b11001011101101:	sigmoid_prime = 18'b000000000101111010;
		14'b11001011101110:	sigmoid_prime = 18'b000000000101111011;
		14'b11001011101111:	sigmoid_prime = 18'b000000000101111100;
		14'b11001011110000:	sigmoid_prime = 18'b000000000101111100;
		14'b11001011110001:	sigmoid_prime = 18'b000000000101111101;
		14'b11001011110010:	sigmoid_prime = 18'b000000000101111110;
		14'b11001011110011:	sigmoid_prime = 18'b000000000101111111;
		14'b11001011110100:	sigmoid_prime = 18'b000000000101111111;
		14'b11001011110101:	sigmoid_prime = 18'b000000000110000000;
		14'b11001011110110:	sigmoid_prime = 18'b000000000110000001;
		14'b11001011110111:	sigmoid_prime = 18'b000000000110000010;
		14'b11001011111000:	sigmoid_prime = 18'b000000000110000010;
		14'b11001011111001:	sigmoid_prime = 18'b000000000110000011;
		14'b11001011111010:	sigmoid_prime = 18'b000000000110000100;
		14'b11001011111011:	sigmoid_prime = 18'b000000000110000101;
		14'b11001011111100:	sigmoid_prime = 18'b000000000110000101;
		14'b11001011111101:	sigmoid_prime = 18'b000000000110000110;
		14'b11001011111110:	sigmoid_prime = 18'b000000000110000111;
		14'b11001011111111:	sigmoid_prime = 18'b000000000110001000;
		14'b11001100000000:	sigmoid_prime = 18'b000000000110001000;
		14'b11001100000001:	sigmoid_prime = 18'b000000000110001001;
		14'b11001100000010:	sigmoid_prime = 18'b000000000110001010;
		14'b11001100000011:	sigmoid_prime = 18'b000000000110001011;
		14'b11001100000100:	sigmoid_prime = 18'b000000000110001100;
		14'b11001100000101:	sigmoid_prime = 18'b000000000110001100;
		14'b11001100000110:	sigmoid_prime = 18'b000000000110001101;
		14'b11001100000111:	sigmoid_prime = 18'b000000000110001110;
		14'b11001100001000:	sigmoid_prime = 18'b000000000110001111;
		14'b11001100001001:	sigmoid_prime = 18'b000000000110001111;
		14'b11001100001010:	sigmoid_prime = 18'b000000000110010000;
		14'b11001100001011:	sigmoid_prime = 18'b000000000110010001;
		14'b11001100001100:	sigmoid_prime = 18'b000000000110010010;
		14'b11001100001101:	sigmoid_prime = 18'b000000000110010011;
		14'b11001100001110:	sigmoid_prime = 18'b000000000110010011;
		14'b11001100001111:	sigmoid_prime = 18'b000000000110010100;
		14'b11001100010000:	sigmoid_prime = 18'b000000000110010101;
		14'b11001100010001:	sigmoid_prime = 18'b000000000110010110;
		14'b11001100010010:	sigmoid_prime = 18'b000000000110010110;
		14'b11001100010011:	sigmoid_prime = 18'b000000000110010111;
		14'b11001100010100:	sigmoid_prime = 18'b000000000110011000;
		14'b11001100010101:	sigmoid_prime = 18'b000000000110011001;
		14'b11001100010110:	sigmoid_prime = 18'b000000000110011010;
		14'b11001100010111:	sigmoid_prime = 18'b000000000110011010;
		14'b11001100011000:	sigmoid_prime = 18'b000000000110011011;
		14'b11001100011001:	sigmoid_prime = 18'b000000000110011100;
		14'b11001100011010:	sigmoid_prime = 18'b000000000110011101;
		14'b11001100011011:	sigmoid_prime = 18'b000000000110011110;
		14'b11001100011100:	sigmoid_prime = 18'b000000000110011110;
		14'b11001100011101:	sigmoid_prime = 18'b000000000110011111;
		14'b11001100011110:	sigmoid_prime = 18'b000000000110100000;
		14'b11001100011111:	sigmoid_prime = 18'b000000000110100001;
		14'b11001100100000:	sigmoid_prime = 18'b000000000110100010;
		14'b11001100100001:	sigmoid_prime = 18'b000000000110100011;
		14'b11001100100010:	sigmoid_prime = 18'b000000000110100011;
		14'b11001100100011:	sigmoid_prime = 18'b000000000110100100;
		14'b11001100100100:	sigmoid_prime = 18'b000000000110100101;
		14'b11001100100101:	sigmoid_prime = 18'b000000000110100110;
		14'b11001100100110:	sigmoid_prime = 18'b000000000110100111;
		14'b11001100100111:	sigmoid_prime = 18'b000000000110100111;
		14'b11001100101000:	sigmoid_prime = 18'b000000000110101000;
		14'b11001100101001:	sigmoid_prime = 18'b000000000110101001;
		14'b11001100101010:	sigmoid_prime = 18'b000000000110101010;
		14'b11001100101011:	sigmoid_prime = 18'b000000000110101011;
		14'b11001100101100:	sigmoid_prime = 18'b000000000110101100;
		14'b11001100101101:	sigmoid_prime = 18'b000000000110101100;
		14'b11001100101110:	sigmoid_prime = 18'b000000000110101101;
		14'b11001100101111:	sigmoid_prime = 18'b000000000110101110;
		14'b11001100110000:	sigmoid_prime = 18'b000000000110101111;
		14'b11001100110001:	sigmoid_prime = 18'b000000000110110000;
		14'b11001100110010:	sigmoid_prime = 18'b000000000110110001;
		14'b11001100110011:	sigmoid_prime = 18'b000000000110110001;
		14'b11001100110100:	sigmoid_prime = 18'b000000000110110010;
		14'b11001100110101:	sigmoid_prime = 18'b000000000110110011;
		14'b11001100110110:	sigmoid_prime = 18'b000000000110110100;
		14'b11001100110111:	sigmoid_prime = 18'b000000000110110101;
		14'b11001100111000:	sigmoid_prime = 18'b000000000110110110;
		14'b11001100111001:	sigmoid_prime = 18'b000000000110110111;
		14'b11001100111010:	sigmoid_prime = 18'b000000000110110111;
		14'b11001100111011:	sigmoid_prime = 18'b000000000110111000;
		14'b11001100111100:	sigmoid_prime = 18'b000000000110111001;
		14'b11001100111101:	sigmoid_prime = 18'b000000000110111010;
		14'b11001100111110:	sigmoid_prime = 18'b000000000110111011;
		14'b11001100111111:	sigmoid_prime = 18'b000000000110111100;
		14'b11001101000000:	sigmoid_prime = 18'b000000000110111101;
		14'b11001101000001:	sigmoid_prime = 18'b000000000110111101;
		14'b11001101000010:	sigmoid_prime = 18'b000000000110111110;
		14'b11001101000011:	sigmoid_prime = 18'b000000000110111111;
		14'b11001101000100:	sigmoid_prime = 18'b000000000111000000;
		14'b11001101000101:	sigmoid_prime = 18'b000000000111000001;
		14'b11001101000110:	sigmoid_prime = 18'b000000000111000010;
		14'b11001101000111:	sigmoid_prime = 18'b000000000111000011;
		14'b11001101001000:	sigmoid_prime = 18'b000000000111000100;
		14'b11001101001001:	sigmoid_prime = 18'b000000000111000100;
		14'b11001101001010:	sigmoid_prime = 18'b000000000111000101;
		14'b11001101001011:	sigmoid_prime = 18'b000000000111000110;
		14'b11001101001100:	sigmoid_prime = 18'b000000000111000111;
		14'b11001101001101:	sigmoid_prime = 18'b000000000111001000;
		14'b11001101001110:	sigmoid_prime = 18'b000000000111001001;
		14'b11001101001111:	sigmoid_prime = 18'b000000000111001010;
		14'b11001101010000:	sigmoid_prime = 18'b000000000111001011;
		14'b11001101010001:	sigmoid_prime = 18'b000000000111001100;
		14'b11001101010010:	sigmoid_prime = 18'b000000000111001100;
		14'b11001101010011:	sigmoid_prime = 18'b000000000111001101;
		14'b11001101010100:	sigmoid_prime = 18'b000000000111001110;
		14'b11001101010101:	sigmoid_prime = 18'b000000000111001111;
		14'b11001101010110:	sigmoid_prime = 18'b000000000111010000;
		14'b11001101010111:	sigmoid_prime = 18'b000000000111010001;
		14'b11001101011000:	sigmoid_prime = 18'b000000000111010010;
		14'b11001101011001:	sigmoid_prime = 18'b000000000111010011;
		14'b11001101011010:	sigmoid_prime = 18'b000000000111010100;
		14'b11001101011011:	sigmoid_prime = 18'b000000000111010101;
		14'b11001101011100:	sigmoid_prime = 18'b000000000111010110;
		14'b11001101011101:	sigmoid_prime = 18'b000000000111010110;
		14'b11001101011110:	sigmoid_prime = 18'b000000000111010111;
		14'b11001101011111:	sigmoid_prime = 18'b000000000111011000;
		14'b11001101100000:	sigmoid_prime = 18'b000000000111011001;
		14'b11001101100001:	sigmoid_prime = 18'b000000000111011010;
		14'b11001101100010:	sigmoid_prime = 18'b000000000111011011;
		14'b11001101100011:	sigmoid_prime = 18'b000000000111011100;
		14'b11001101100100:	sigmoid_prime = 18'b000000000111011101;
		14'b11001101100101:	sigmoid_prime = 18'b000000000111011110;
		14'b11001101100110:	sigmoid_prime = 18'b000000000111011111;
		14'b11001101100111:	sigmoid_prime = 18'b000000000111100000;
		14'b11001101101000:	sigmoid_prime = 18'b000000000111100001;
		14'b11001101101001:	sigmoid_prime = 18'b000000000111100010;
		14'b11001101101010:	sigmoid_prime = 18'b000000000111100010;
		14'b11001101101011:	sigmoid_prime = 18'b000000000111100011;
		14'b11001101101100:	sigmoid_prime = 18'b000000000111100100;
		14'b11001101101101:	sigmoid_prime = 18'b000000000111100101;
		14'b11001101101110:	sigmoid_prime = 18'b000000000111100110;
		14'b11001101101111:	sigmoid_prime = 18'b000000000111100111;
		14'b11001101110000:	sigmoid_prime = 18'b000000000111101000;
		14'b11001101110001:	sigmoid_prime = 18'b000000000111101001;
		14'b11001101110010:	sigmoid_prime = 18'b000000000111101010;
		14'b11001101110011:	sigmoid_prime = 18'b000000000111101011;
		14'b11001101110100:	sigmoid_prime = 18'b000000000111101100;
		14'b11001101110101:	sigmoid_prime = 18'b000000000111101101;
		14'b11001101110110:	sigmoid_prime = 18'b000000000111101110;
		14'b11001101110111:	sigmoid_prime = 18'b000000000111101111;
		14'b11001101111000:	sigmoid_prime = 18'b000000000111110000;
		14'b11001101111001:	sigmoid_prime = 18'b000000000111110001;
		14'b11001101111010:	sigmoid_prime = 18'b000000000111110010;
		14'b11001101111011:	sigmoid_prime = 18'b000000000111110011;
		14'b11001101111100:	sigmoid_prime = 18'b000000000111110100;
		14'b11001101111101:	sigmoid_prime = 18'b000000000111110101;
		14'b11001101111110:	sigmoid_prime = 18'b000000000111110110;
		14'b11001101111111:	sigmoid_prime = 18'b000000000111110111;
		14'b11001110000000:	sigmoid_prime = 18'b000000000111111000;
		14'b11001110000001:	sigmoid_prime = 18'b000000000111111001;
		14'b11001110000010:	sigmoid_prime = 18'b000000000111111010;
		14'b11001110000011:	sigmoid_prime = 18'b000000000111111011;
		14'b11001110000100:	sigmoid_prime = 18'b000000000111111100;
		14'b11001110000101:	sigmoid_prime = 18'b000000000111111101;
		14'b11001110000110:	sigmoid_prime = 18'b000000000111111110;
		14'b11001110000111:	sigmoid_prime = 18'b000000000111111111;
		14'b11001110001000:	sigmoid_prime = 18'b000000001000000000;
		14'b11001110001001:	sigmoid_prime = 18'b000000001000000001;
		14'b11001110001010:	sigmoid_prime = 18'b000000001000000010;
		14'b11001110001011:	sigmoid_prime = 18'b000000001000000011;
		14'b11001110001100:	sigmoid_prime = 18'b000000001000000100;
		14'b11001110001101:	sigmoid_prime = 18'b000000001000000101;
		14'b11001110001110:	sigmoid_prime = 18'b000000001000000110;
		14'b11001110001111:	sigmoid_prime = 18'b000000001000000111;
		14'b11001110010000:	sigmoid_prime = 18'b000000001000001000;
		14'b11001110010001:	sigmoid_prime = 18'b000000001000001001;
		14'b11001110010010:	sigmoid_prime = 18'b000000001000001010;
		14'b11001110010011:	sigmoid_prime = 18'b000000001000001011;
		14'b11001110010100:	sigmoid_prime = 18'b000000001000001100;
		14'b11001110010101:	sigmoid_prime = 18'b000000001000001101;
		14'b11001110010110:	sigmoid_prime = 18'b000000001000001110;
		14'b11001110010111:	sigmoid_prime = 18'b000000001000001111;
		14'b11001110011000:	sigmoid_prime = 18'b000000001000010000;
		14'b11001110011001:	sigmoid_prime = 18'b000000001000010001;
		14'b11001110011010:	sigmoid_prime = 18'b000000001000010010;
		14'b11001110011011:	sigmoid_prime = 18'b000000001000010011;
		14'b11001110011100:	sigmoid_prime = 18'b000000001000010100;
		14'b11001110011101:	sigmoid_prime = 18'b000000001000010101;
		14'b11001110011110:	sigmoid_prime = 18'b000000001000010110;
		14'b11001110011111:	sigmoid_prime = 18'b000000001000010111;
		14'b11001110100000:	sigmoid_prime = 18'b000000001000011000;
		14'b11001110100001:	sigmoid_prime = 18'b000000001000011001;
		14'b11001110100010:	sigmoid_prime = 18'b000000001000011010;
		14'b11001110100011:	sigmoid_prime = 18'b000000001000011011;
		14'b11001110100100:	sigmoid_prime = 18'b000000001000011100;
		14'b11001110100101:	sigmoid_prime = 18'b000000001000011101;
		14'b11001110100110:	sigmoid_prime = 18'b000000001000011110;
		14'b11001110100111:	sigmoid_prime = 18'b000000001000011111;
		14'b11001110101000:	sigmoid_prime = 18'b000000001000100000;
		14'b11001110101001:	sigmoid_prime = 18'b000000001000100001;
		14'b11001110101010:	sigmoid_prime = 18'b000000001000100011;
		14'b11001110101011:	sigmoid_prime = 18'b000000001000100100;
		14'b11001110101100:	sigmoid_prime = 18'b000000001000100101;
		14'b11001110101101:	sigmoid_prime = 18'b000000001000100110;
		14'b11001110101110:	sigmoid_prime = 18'b000000001000100111;
		14'b11001110101111:	sigmoid_prime = 18'b000000001000101000;
		14'b11001110110000:	sigmoid_prime = 18'b000000001000101001;
		14'b11001110110001:	sigmoid_prime = 18'b000000001000101010;
		14'b11001110110010:	sigmoid_prime = 18'b000000001000101011;
		14'b11001110110011:	sigmoid_prime = 18'b000000001000101100;
		14'b11001110110100:	sigmoid_prime = 18'b000000001000101101;
		14'b11001110110101:	sigmoid_prime = 18'b000000001000101110;
		14'b11001110110110:	sigmoid_prime = 18'b000000001000101111;
		14'b11001110110111:	sigmoid_prime = 18'b000000001000110001;
		14'b11001110111000:	sigmoid_prime = 18'b000000001000110010;
		14'b11001110111001:	sigmoid_prime = 18'b000000001000110011;
		14'b11001110111010:	sigmoid_prime = 18'b000000001000110100;
		14'b11001110111011:	sigmoid_prime = 18'b000000001000110101;
		14'b11001110111100:	sigmoid_prime = 18'b000000001000110110;
		14'b11001110111101:	sigmoid_prime = 18'b000000001000110111;
		14'b11001110111110:	sigmoid_prime = 18'b000000001000111000;
		14'b11001110111111:	sigmoid_prime = 18'b000000001000111001;
		14'b11001111000000:	sigmoid_prime = 18'b000000001000111010;
		14'b11001111000001:	sigmoid_prime = 18'b000000001000111100;
		14'b11001111000010:	sigmoid_prime = 18'b000000001000111101;
		14'b11001111000011:	sigmoid_prime = 18'b000000001000111110;
		14'b11001111000100:	sigmoid_prime = 18'b000000001000111111;
		14'b11001111000101:	sigmoid_prime = 18'b000000001001000000;
		14'b11001111000110:	sigmoid_prime = 18'b000000001001000001;
		14'b11001111000111:	sigmoid_prime = 18'b000000001001000010;
		14'b11001111001000:	sigmoid_prime = 18'b000000001001000011;
		14'b11001111001001:	sigmoid_prime = 18'b000000001001000101;
		14'b11001111001010:	sigmoid_prime = 18'b000000001001000110;
		14'b11001111001011:	sigmoid_prime = 18'b000000001001000111;
		14'b11001111001100:	sigmoid_prime = 18'b000000001001001000;
		14'b11001111001101:	sigmoid_prime = 18'b000000001001001001;
		14'b11001111001110:	sigmoid_prime = 18'b000000001001001010;
		14'b11001111001111:	sigmoid_prime = 18'b000000001001001011;
		14'b11001111010000:	sigmoid_prime = 18'b000000001001001100;
		14'b11001111010001:	sigmoid_prime = 18'b000000001001001110;
		14'b11001111010010:	sigmoid_prime = 18'b000000001001001111;
		14'b11001111010011:	sigmoid_prime = 18'b000000001001010000;
		14'b11001111010100:	sigmoid_prime = 18'b000000001001010001;
		14'b11001111010101:	sigmoid_prime = 18'b000000001001010010;
		14'b11001111010110:	sigmoid_prime = 18'b000000001001010011;
		14'b11001111010111:	sigmoid_prime = 18'b000000001001010101;
		14'b11001111011000:	sigmoid_prime = 18'b000000001001010110;
		14'b11001111011001:	sigmoid_prime = 18'b000000001001010111;
		14'b11001111011010:	sigmoid_prime = 18'b000000001001011000;
		14'b11001111011011:	sigmoid_prime = 18'b000000001001011001;
		14'b11001111011100:	sigmoid_prime = 18'b000000001001011010;
		14'b11001111011101:	sigmoid_prime = 18'b000000001001011100;
		14'b11001111011110:	sigmoid_prime = 18'b000000001001011101;
		14'b11001111011111:	sigmoid_prime = 18'b000000001001011110;
		14'b11001111100000:	sigmoid_prime = 18'b000000001001011111;
		14'b11001111100001:	sigmoid_prime = 18'b000000001001100000;
		14'b11001111100010:	sigmoid_prime = 18'b000000001001100001;
		14'b11001111100011:	sigmoid_prime = 18'b000000001001100011;
		14'b11001111100100:	sigmoid_prime = 18'b000000001001100100;
		14'b11001111100101:	sigmoid_prime = 18'b000000001001100101;
		14'b11001111100110:	sigmoid_prime = 18'b000000001001100110;
		14'b11001111100111:	sigmoid_prime = 18'b000000001001100111;
		14'b11001111101000:	sigmoid_prime = 18'b000000001001101001;
		14'b11001111101001:	sigmoid_prime = 18'b000000001001101010;
		14'b11001111101010:	sigmoid_prime = 18'b000000001001101011;
		14'b11001111101011:	sigmoid_prime = 18'b000000001001101100;
		14'b11001111101100:	sigmoid_prime = 18'b000000001001101101;
		14'b11001111101101:	sigmoid_prime = 18'b000000001001101111;
		14'b11001111101110:	sigmoid_prime = 18'b000000001001110000;
		14'b11001111101111:	sigmoid_prime = 18'b000000001001110001;
		14'b11001111110000:	sigmoid_prime = 18'b000000001001110010;
		14'b11001111110001:	sigmoid_prime = 18'b000000001001110100;
		14'b11001111110010:	sigmoid_prime = 18'b000000001001110101;
		14'b11001111110011:	sigmoid_prime = 18'b000000001001110110;
		14'b11001111110100:	sigmoid_prime = 18'b000000001001110111;
		14'b11001111110101:	sigmoid_prime = 18'b000000001001111000;
		14'b11001111110110:	sigmoid_prime = 18'b000000001001111010;
		14'b11001111110111:	sigmoid_prime = 18'b000000001001111011;
		14'b11001111111000:	sigmoid_prime = 18'b000000001001111100;
		14'b11001111111001:	sigmoid_prime = 18'b000000001001111101;
		14'b11001111111010:	sigmoid_prime = 18'b000000001001111111;
		14'b11001111111011:	sigmoid_prime = 18'b000000001010000000;
		14'b11001111111100:	sigmoid_prime = 18'b000000001010000001;
		14'b11001111111101:	sigmoid_prime = 18'b000000001010000010;
		14'b11001111111110:	sigmoid_prime = 18'b000000001010000100;
		14'b11001111111111:	sigmoid_prime = 18'b000000001010000101;
		14'b11010000000000:	sigmoid_prime = 18'b000000001010000110;
		14'b11010000000001:	sigmoid_prime = 18'b000000001010000111;
		14'b11010000000010:	sigmoid_prime = 18'b000000001010001001;
		14'b11010000000011:	sigmoid_prime = 18'b000000001010001010;
		14'b11010000000100:	sigmoid_prime = 18'b000000001010001011;
		14'b11010000000101:	sigmoid_prime = 18'b000000001010001100;
		14'b11010000000110:	sigmoid_prime = 18'b000000001010001110;
		14'b11010000000111:	sigmoid_prime = 18'b000000001010001111;
		14'b11010000001000:	sigmoid_prime = 18'b000000001010010000;
		14'b11010000001001:	sigmoid_prime = 18'b000000001010010001;
		14'b11010000001010:	sigmoid_prime = 18'b000000001010010011;
		14'b11010000001011:	sigmoid_prime = 18'b000000001010010100;
		14'b11010000001100:	sigmoid_prime = 18'b000000001010010101;
		14'b11010000001101:	sigmoid_prime = 18'b000000001010010111;
		14'b11010000001110:	sigmoid_prime = 18'b000000001010011000;
		14'b11010000001111:	sigmoid_prime = 18'b000000001010011001;
		14'b11010000010000:	sigmoid_prime = 18'b000000001010011011;
		14'b11010000010001:	sigmoid_prime = 18'b000000001010011100;
		14'b11010000010010:	sigmoid_prime = 18'b000000001010011101;
		14'b11010000010011:	sigmoid_prime = 18'b000000001010011110;
		14'b11010000010100:	sigmoid_prime = 18'b000000001010100000;
		14'b11010000010101:	sigmoid_prime = 18'b000000001010100001;
		14'b11010000010110:	sigmoid_prime = 18'b000000001010100010;
		14'b11010000010111:	sigmoid_prime = 18'b000000001010100100;
		14'b11010000011000:	sigmoid_prime = 18'b000000001010100101;
		14'b11010000011001:	sigmoid_prime = 18'b000000001010100110;
		14'b11010000011010:	sigmoid_prime = 18'b000000001010101000;
		14'b11010000011011:	sigmoid_prime = 18'b000000001010101001;
		14'b11010000011100:	sigmoid_prime = 18'b000000001010101010;
		14'b11010000011101:	sigmoid_prime = 18'b000000001010101100;
		14'b11010000011110:	sigmoid_prime = 18'b000000001010101101;
		14'b11010000011111:	sigmoid_prime = 18'b000000001010101110;
		14'b11010000100000:	sigmoid_prime = 18'b000000001010110000;
		14'b11010000100001:	sigmoid_prime = 18'b000000001010110001;
		14'b11010000100010:	sigmoid_prime = 18'b000000001010110010;
		14'b11010000100011:	sigmoid_prime = 18'b000000001010110100;
		14'b11010000100100:	sigmoid_prime = 18'b000000001010110101;
		14'b11010000100101:	sigmoid_prime = 18'b000000001010110110;
		14'b11010000100110:	sigmoid_prime = 18'b000000001010111000;
		14'b11010000100111:	sigmoid_prime = 18'b000000001010111001;
		14'b11010000101000:	sigmoid_prime = 18'b000000001010111010;
		14'b11010000101001:	sigmoid_prime = 18'b000000001010111100;
		14'b11010000101010:	sigmoid_prime = 18'b000000001010111101;
		14'b11010000101011:	sigmoid_prime = 18'b000000001010111110;
		14'b11010000101100:	sigmoid_prime = 18'b000000001011000000;
		14'b11010000101101:	sigmoid_prime = 18'b000000001011000001;
		14'b11010000101110:	sigmoid_prime = 18'b000000001011000011;
		14'b11010000101111:	sigmoid_prime = 18'b000000001011000100;
		14'b11010000110000:	sigmoid_prime = 18'b000000001011000101;
		14'b11010000110001:	sigmoid_prime = 18'b000000001011000111;
		14'b11010000110010:	sigmoid_prime = 18'b000000001011001000;
		14'b11010000110011:	sigmoid_prime = 18'b000000001011001001;
		14'b11010000110100:	sigmoid_prime = 18'b000000001011001011;
		14'b11010000110101:	sigmoid_prime = 18'b000000001011001100;
		14'b11010000110110:	sigmoid_prime = 18'b000000001011001110;
		14'b11010000110111:	sigmoid_prime = 18'b000000001011001111;
		14'b11010000111000:	sigmoid_prime = 18'b000000001011010000;
		14'b11010000111001:	sigmoid_prime = 18'b000000001011010010;
		14'b11010000111010:	sigmoid_prime = 18'b000000001011010011;
		14'b11010000111011:	sigmoid_prime = 18'b000000001011010101;
		14'b11010000111100:	sigmoid_prime = 18'b000000001011010110;
		14'b11010000111101:	sigmoid_prime = 18'b000000001011010111;
		14'b11010000111110:	sigmoid_prime = 18'b000000001011011001;
		14'b11010000111111:	sigmoid_prime = 18'b000000001011011010;
		14'b11010001000000:	sigmoid_prime = 18'b000000001011011100;
		14'b11010001000001:	sigmoid_prime = 18'b000000001011011101;
		14'b11010001000010:	sigmoid_prime = 18'b000000001011011111;
		14'b11010001000011:	sigmoid_prime = 18'b000000001011100000;
		14'b11010001000100:	sigmoid_prime = 18'b000000001011100001;
		14'b11010001000101:	sigmoid_prime = 18'b000000001011100011;
		14'b11010001000110:	sigmoid_prime = 18'b000000001011100100;
		14'b11010001000111:	sigmoid_prime = 18'b000000001011100110;
		14'b11010001001000:	sigmoid_prime = 18'b000000001011100111;
		14'b11010001001001:	sigmoid_prime = 18'b000000001011101001;
		14'b11010001001010:	sigmoid_prime = 18'b000000001011101010;
		14'b11010001001011:	sigmoid_prime = 18'b000000001011101011;
		14'b11010001001100:	sigmoid_prime = 18'b000000001011101101;
		14'b11010001001101:	sigmoid_prime = 18'b000000001011101110;
		14'b11010001001110:	sigmoid_prime = 18'b000000001011110000;
		14'b11010001001111:	sigmoid_prime = 18'b000000001011110001;
		14'b11010001010000:	sigmoid_prime = 18'b000000001011110011;
		14'b11010001010001:	sigmoid_prime = 18'b000000001011110100;
		14'b11010001010010:	sigmoid_prime = 18'b000000001011110110;
		14'b11010001010011:	sigmoid_prime = 18'b000000001011110111;
		14'b11010001010100:	sigmoid_prime = 18'b000000001011111001;
		14'b11010001010101:	sigmoid_prime = 18'b000000001011111010;
		14'b11010001010110:	sigmoid_prime = 18'b000000001011111100;
		14'b11010001010111:	sigmoid_prime = 18'b000000001011111101;
		14'b11010001011000:	sigmoid_prime = 18'b000000001011111111;
		14'b11010001011001:	sigmoid_prime = 18'b000000001100000000;
		14'b11010001011010:	sigmoid_prime = 18'b000000001100000010;
		14'b11010001011011:	sigmoid_prime = 18'b000000001100000011;
		14'b11010001011100:	sigmoid_prime = 18'b000000001100000101;
		14'b11010001011101:	sigmoid_prime = 18'b000000001100000110;
		14'b11010001011110:	sigmoid_prime = 18'b000000001100001000;
		14'b11010001011111:	sigmoid_prime = 18'b000000001100001001;
		14'b11010001100000:	sigmoid_prime = 18'b000000001100001011;
		14'b11010001100001:	sigmoid_prime = 18'b000000001100001100;
		14'b11010001100010:	sigmoid_prime = 18'b000000001100001110;
		14'b11010001100011:	sigmoid_prime = 18'b000000001100001111;
		14'b11010001100100:	sigmoid_prime = 18'b000000001100010001;
		14'b11010001100101:	sigmoid_prime = 18'b000000001100010010;
		14'b11010001100110:	sigmoid_prime = 18'b000000001100010100;
		14'b11010001100111:	sigmoid_prime = 18'b000000001100010101;
		14'b11010001101000:	sigmoid_prime = 18'b000000001100010111;
		14'b11010001101001:	sigmoid_prime = 18'b000000001100011000;
		14'b11010001101010:	sigmoid_prime = 18'b000000001100011010;
		14'b11010001101011:	sigmoid_prime = 18'b000000001100011011;
		14'b11010001101100:	sigmoid_prime = 18'b000000001100011101;
		14'b11010001101101:	sigmoid_prime = 18'b000000001100011111;
		14'b11010001101110:	sigmoid_prime = 18'b000000001100100000;
		14'b11010001101111:	sigmoid_prime = 18'b000000001100100010;
		14'b11010001110000:	sigmoid_prime = 18'b000000001100100011;
		14'b11010001110001:	sigmoid_prime = 18'b000000001100100101;
		14'b11010001110010:	sigmoid_prime = 18'b000000001100100110;
		14'b11010001110011:	sigmoid_prime = 18'b000000001100101000;
		14'b11010001110100:	sigmoid_prime = 18'b000000001100101001;
		14'b11010001110101:	sigmoid_prime = 18'b000000001100101011;
		14'b11010001110110:	sigmoid_prime = 18'b000000001100101101;
		14'b11010001110111:	sigmoid_prime = 18'b000000001100101110;
		14'b11010001111000:	sigmoid_prime = 18'b000000001100110000;
		14'b11010001111001:	sigmoid_prime = 18'b000000001100110001;
		14'b11010001111010:	sigmoid_prime = 18'b000000001100110011;
		14'b11010001111011:	sigmoid_prime = 18'b000000001100110101;
		14'b11010001111100:	sigmoid_prime = 18'b000000001100110110;
		14'b11010001111101:	sigmoid_prime = 18'b000000001100111000;
		14'b11010001111110:	sigmoid_prime = 18'b000000001100111001;
		14'b11010001111111:	sigmoid_prime = 18'b000000001100111011;
		14'b11010010000000:	sigmoid_prime = 18'b000000001100111101;
		14'b11010010000001:	sigmoid_prime = 18'b000000001100111110;
		14'b11010010000010:	sigmoid_prime = 18'b000000001101000000;
		14'b11010010000011:	sigmoid_prime = 18'b000000001101000001;
		14'b11010010000100:	sigmoid_prime = 18'b000000001101000011;
		14'b11010010000101:	sigmoid_prime = 18'b000000001101000101;
		14'b11010010000110:	sigmoid_prime = 18'b000000001101000110;
		14'b11010010000111:	sigmoid_prime = 18'b000000001101001000;
		14'b11010010001000:	sigmoid_prime = 18'b000000001101001010;
		14'b11010010001001:	sigmoid_prime = 18'b000000001101001011;
		14'b11010010001010:	sigmoid_prime = 18'b000000001101001101;
		14'b11010010001011:	sigmoid_prime = 18'b000000001101001110;
		14'b11010010001100:	sigmoid_prime = 18'b000000001101010000;
		14'b11010010001101:	sigmoid_prime = 18'b000000001101010010;
		14'b11010010001110:	sigmoid_prime = 18'b000000001101010011;
		14'b11010010001111:	sigmoid_prime = 18'b000000001101010101;
		14'b11010010010000:	sigmoid_prime = 18'b000000001101010111;
		14'b11010010010001:	sigmoid_prime = 18'b000000001101011000;
		14'b11010010010010:	sigmoid_prime = 18'b000000001101011010;
		14'b11010010010011:	sigmoid_prime = 18'b000000001101011100;
		14'b11010010010100:	sigmoid_prime = 18'b000000001101011101;
		14'b11010010010101:	sigmoid_prime = 18'b000000001101011111;
		14'b11010010010110:	sigmoid_prime = 18'b000000001101100001;
		14'b11010010010111:	sigmoid_prime = 18'b000000001101100010;
		14'b11010010011000:	sigmoid_prime = 18'b000000001101100100;
		14'b11010010011001:	sigmoid_prime = 18'b000000001101100110;
		14'b11010010011010:	sigmoid_prime = 18'b000000001101100111;
		14'b11010010011011:	sigmoid_prime = 18'b000000001101101001;
		14'b11010010011100:	sigmoid_prime = 18'b000000001101101011;
		14'b11010010011101:	sigmoid_prime = 18'b000000001101101101;
		14'b11010010011110:	sigmoid_prime = 18'b000000001101101110;
		14'b11010010011111:	sigmoid_prime = 18'b000000001101110000;
		14'b11010010100000:	sigmoid_prime = 18'b000000001101110010;
		14'b11010010100001:	sigmoid_prime = 18'b000000001101110011;
		14'b11010010100010:	sigmoid_prime = 18'b000000001101110101;
		14'b11010010100011:	sigmoid_prime = 18'b000000001101110111;
		14'b11010010100100:	sigmoid_prime = 18'b000000001101111001;
		14'b11010010100101:	sigmoid_prime = 18'b000000001101111010;
		14'b11010010100110:	sigmoid_prime = 18'b000000001101111100;
		14'b11010010100111:	sigmoid_prime = 18'b000000001101111110;
		14'b11010010101000:	sigmoid_prime = 18'b000000001101111111;
		14'b11010010101001:	sigmoid_prime = 18'b000000001110000001;
		14'b11010010101010:	sigmoid_prime = 18'b000000001110000011;
		14'b11010010101011:	sigmoid_prime = 18'b000000001110000101;
		14'b11010010101100:	sigmoid_prime = 18'b000000001110000110;
		14'b11010010101101:	sigmoid_prime = 18'b000000001110001000;
		14'b11010010101110:	sigmoid_prime = 18'b000000001110001010;
		14'b11010010101111:	sigmoid_prime = 18'b000000001110001100;
		14'b11010010110000:	sigmoid_prime = 18'b000000001110001101;
		14'b11010010110001:	sigmoid_prime = 18'b000000001110001111;
		14'b11010010110010:	sigmoid_prime = 18'b000000001110010001;
		14'b11010010110011:	sigmoid_prime = 18'b000000001110010011;
		14'b11010010110100:	sigmoid_prime = 18'b000000001110010101;
		14'b11010010110101:	sigmoid_prime = 18'b000000001110010110;
		14'b11010010110110:	sigmoid_prime = 18'b000000001110011000;
		14'b11010010110111:	sigmoid_prime = 18'b000000001110011010;
		14'b11010010111000:	sigmoid_prime = 18'b000000001110011100;
		14'b11010010111001:	sigmoid_prime = 18'b000000001110011110;
		14'b11010010111010:	sigmoid_prime = 18'b000000001110011111;
		14'b11010010111011:	sigmoid_prime = 18'b000000001110100001;
		14'b11010010111100:	sigmoid_prime = 18'b000000001110100011;
		14'b11010010111101:	sigmoid_prime = 18'b000000001110100101;
		14'b11010010111110:	sigmoid_prime = 18'b000000001110100111;
		14'b11010010111111:	sigmoid_prime = 18'b000000001110101000;
		14'b11010011000000:	sigmoid_prime = 18'b000000001110101010;
		14'b11010011000001:	sigmoid_prime = 18'b000000001110101100;
		14'b11010011000010:	sigmoid_prime = 18'b000000001110101110;
		14'b11010011000011:	sigmoid_prime = 18'b000000001110110000;
		14'b11010011000100:	sigmoid_prime = 18'b000000001110110001;
		14'b11010011000101:	sigmoid_prime = 18'b000000001110110011;
		14'b11010011000110:	sigmoid_prime = 18'b000000001110110101;
		14'b11010011000111:	sigmoid_prime = 18'b000000001110110111;
		14'b11010011001000:	sigmoid_prime = 18'b000000001110111001;
		14'b11010011001001:	sigmoid_prime = 18'b000000001110111011;
		14'b11010011001010:	sigmoid_prime = 18'b000000001110111101;
		14'b11010011001011:	sigmoid_prime = 18'b000000001110111110;
		14'b11010011001100:	sigmoid_prime = 18'b000000001111000000;
		14'b11010011001101:	sigmoid_prime = 18'b000000001111000010;
		14'b11010011001110:	sigmoid_prime = 18'b000000001111000100;
		14'b11010011001111:	sigmoid_prime = 18'b000000001111000110;
		14'b11010011010000:	sigmoid_prime = 18'b000000001111001000;
		14'b11010011010001:	sigmoid_prime = 18'b000000001111001010;
		14'b11010011010010:	sigmoid_prime = 18'b000000001111001011;
		14'b11010011010011:	sigmoid_prime = 18'b000000001111001101;
		14'b11010011010100:	sigmoid_prime = 18'b000000001111001111;
		14'b11010011010101:	sigmoid_prime = 18'b000000001111010001;
		14'b11010011010110:	sigmoid_prime = 18'b000000001111010011;
		14'b11010011010111:	sigmoid_prime = 18'b000000001111010101;
		14'b11010011011000:	sigmoid_prime = 18'b000000001111010111;
		14'b11010011011001:	sigmoid_prime = 18'b000000001111011001;
		14'b11010011011010:	sigmoid_prime = 18'b000000001111011011;
		14'b11010011011011:	sigmoid_prime = 18'b000000001111011101;
		14'b11010011011100:	sigmoid_prime = 18'b000000001111011111;
		14'b11010011011101:	sigmoid_prime = 18'b000000001111100000;
		14'b11010011011110:	sigmoid_prime = 18'b000000001111100010;
		14'b11010011011111:	sigmoid_prime = 18'b000000001111100100;
		14'b11010011100000:	sigmoid_prime = 18'b000000001111100110;
		14'b11010011100001:	sigmoid_prime = 18'b000000001111101000;
		14'b11010011100010:	sigmoid_prime = 18'b000000001111101010;
		14'b11010011100011:	sigmoid_prime = 18'b000000001111101100;
		14'b11010011100100:	sigmoid_prime = 18'b000000001111101110;
		14'b11010011100101:	sigmoid_prime = 18'b000000001111110000;
		14'b11010011100110:	sigmoid_prime = 18'b000000001111110010;
		14'b11010011100111:	sigmoid_prime = 18'b000000001111110100;
		14'b11010011101000:	sigmoid_prime = 18'b000000001111110110;
		14'b11010011101001:	sigmoid_prime = 18'b000000001111111000;
		14'b11010011101010:	sigmoid_prime = 18'b000000001111111010;
		14'b11010011101011:	sigmoid_prime = 18'b000000001111111100;
		14'b11010011101100:	sigmoid_prime = 18'b000000001111111110;
		14'b11010011101101:	sigmoid_prime = 18'b000000010000000000;
		14'b11010011101110:	sigmoid_prime = 18'b000000010000000010;
		14'b11010011101111:	sigmoid_prime = 18'b000000010000000100;
		14'b11010011110000:	sigmoid_prime = 18'b000000010000000110;
		14'b11010011110001:	sigmoid_prime = 18'b000000010000001000;
		14'b11010011110010:	sigmoid_prime = 18'b000000010000001010;
		14'b11010011110011:	sigmoid_prime = 18'b000000010000001100;
		14'b11010011110100:	sigmoid_prime = 18'b000000010000001110;
		14'b11010011110101:	sigmoid_prime = 18'b000000010000010000;
		14'b11010011110110:	sigmoid_prime = 18'b000000010000010010;
		14'b11010011110111:	sigmoid_prime = 18'b000000010000010100;
		14'b11010011111000:	sigmoid_prime = 18'b000000010000010110;
		14'b11010011111001:	sigmoid_prime = 18'b000000010000011000;
		14'b11010011111010:	sigmoid_prime = 18'b000000010000011010;
		14'b11010011111011:	sigmoid_prime = 18'b000000010000011100;
		14'b11010011111100:	sigmoid_prime = 18'b000000010000011110;
		14'b11010011111101:	sigmoid_prime = 18'b000000010000100000;
		14'b11010011111110:	sigmoid_prime = 18'b000000010000100010;
		14'b11010011111111:	sigmoid_prime = 18'b000000010000100100;
		14'b11010100000000:	sigmoid_prime = 18'b000000010000100110;
		14'b11010100000001:	sigmoid_prime = 18'b000000010000101000;
		14'b11010100000010:	sigmoid_prime = 18'b000000010000101010;
		14'b11010100000011:	sigmoid_prime = 18'b000000010000101100;
		14'b11010100000100:	sigmoid_prime = 18'b000000010000101110;
		14'b11010100000101:	sigmoid_prime = 18'b000000010000110000;
		14'b11010100000110:	sigmoid_prime = 18'b000000010000110011;
		14'b11010100000111:	sigmoid_prime = 18'b000000010000110101;
		14'b11010100001000:	sigmoid_prime = 18'b000000010000110111;
		14'b11010100001001:	sigmoid_prime = 18'b000000010000111001;
		14'b11010100001010:	sigmoid_prime = 18'b000000010000111011;
		14'b11010100001011:	sigmoid_prime = 18'b000000010000111101;
		14'b11010100001100:	sigmoid_prime = 18'b000000010000111111;
		14'b11010100001101:	sigmoid_prime = 18'b000000010001000001;
		14'b11010100001110:	sigmoid_prime = 18'b000000010001000011;
		14'b11010100001111:	sigmoid_prime = 18'b000000010001000101;
		14'b11010100010000:	sigmoid_prime = 18'b000000010001001000;
		14'b11010100010001:	sigmoid_prime = 18'b000000010001001010;
		14'b11010100010010:	sigmoid_prime = 18'b000000010001001100;
		14'b11010100010011:	sigmoid_prime = 18'b000000010001001110;
		14'b11010100010100:	sigmoid_prime = 18'b000000010001010000;
		14'b11010100010101:	sigmoid_prime = 18'b000000010001010010;
		14'b11010100010110:	sigmoid_prime = 18'b000000010001010100;
		14'b11010100010111:	sigmoid_prime = 18'b000000010001010111;
		14'b11010100011000:	sigmoid_prime = 18'b000000010001011001;
		14'b11010100011001:	sigmoid_prime = 18'b000000010001011011;
		14'b11010100011010:	sigmoid_prime = 18'b000000010001011101;
		14'b11010100011011:	sigmoid_prime = 18'b000000010001011111;
		14'b11010100011100:	sigmoid_prime = 18'b000000010001100001;
		14'b11010100011101:	sigmoid_prime = 18'b000000010001100100;
		14'b11010100011110:	sigmoid_prime = 18'b000000010001100110;
		14'b11010100011111:	sigmoid_prime = 18'b000000010001101000;
		14'b11010100100000:	sigmoid_prime = 18'b000000010001101010;
		14'b11010100100001:	sigmoid_prime = 18'b000000010001101100;
		14'b11010100100010:	sigmoid_prime = 18'b000000010001101110;
		14'b11010100100011:	sigmoid_prime = 18'b000000010001110001;
		14'b11010100100100:	sigmoid_prime = 18'b000000010001110011;
		14'b11010100100101:	sigmoid_prime = 18'b000000010001110101;
		14'b11010100100110:	sigmoid_prime = 18'b000000010001110111;
		14'b11010100100111:	sigmoid_prime = 18'b000000010001111001;
		14'b11010100101000:	sigmoid_prime = 18'b000000010001111100;
		14'b11010100101001:	sigmoid_prime = 18'b000000010001111110;
		14'b11010100101010:	sigmoid_prime = 18'b000000010010000000;
		14'b11010100101011:	sigmoid_prime = 18'b000000010010000010;
		14'b11010100101100:	sigmoid_prime = 18'b000000010010000101;
		14'b11010100101101:	sigmoid_prime = 18'b000000010010000111;
		14'b11010100101110:	sigmoid_prime = 18'b000000010010001001;
		14'b11010100101111:	sigmoid_prime = 18'b000000010010001011;
		14'b11010100110000:	sigmoid_prime = 18'b000000010010001110;
		14'b11010100110001:	sigmoid_prime = 18'b000000010010010000;
		14'b11010100110010:	sigmoid_prime = 18'b000000010010010010;
		14'b11010100110011:	sigmoid_prime = 18'b000000010010010100;
		14'b11010100110100:	sigmoid_prime = 18'b000000010010010111;
		14'b11010100110101:	sigmoid_prime = 18'b000000010010011001;
		14'b11010100110110:	sigmoid_prime = 18'b000000010010011011;
		14'b11010100110111:	sigmoid_prime = 18'b000000010010011110;
		14'b11010100111000:	sigmoid_prime = 18'b000000010010100000;
		14'b11010100111001:	sigmoid_prime = 18'b000000010010100010;
		14'b11010100111010:	sigmoid_prime = 18'b000000010010100100;
		14'b11010100111011:	sigmoid_prime = 18'b000000010010100111;
		14'b11010100111100:	sigmoid_prime = 18'b000000010010101001;
		14'b11010100111101:	sigmoid_prime = 18'b000000010010101011;
		14'b11010100111110:	sigmoid_prime = 18'b000000010010101110;
		14'b11010100111111:	sigmoid_prime = 18'b000000010010110000;
		14'b11010101000000:	sigmoid_prime = 18'b000000010010110010;
		14'b11010101000001:	sigmoid_prime = 18'b000000010010110101;
		14'b11010101000010:	sigmoid_prime = 18'b000000010010110111;
		14'b11010101000011:	sigmoid_prime = 18'b000000010010111001;
		14'b11010101000100:	sigmoid_prime = 18'b000000010010111100;
		14'b11010101000101:	sigmoid_prime = 18'b000000010010111110;
		14'b11010101000110:	sigmoid_prime = 18'b000000010011000000;
		14'b11010101000111:	sigmoid_prime = 18'b000000010011000011;
		14'b11010101001000:	sigmoid_prime = 18'b000000010011000101;
		14'b11010101001001:	sigmoid_prime = 18'b000000010011000111;
		14'b11010101001010:	sigmoid_prime = 18'b000000010011001010;
		14'b11010101001011:	sigmoid_prime = 18'b000000010011001100;
		14'b11010101001100:	sigmoid_prime = 18'b000000010011001111;
		14'b11010101001101:	sigmoid_prime = 18'b000000010011010001;
		14'b11010101001110:	sigmoid_prime = 18'b000000010011010011;
		14'b11010101001111:	sigmoid_prime = 18'b000000010011010110;
		14'b11010101010000:	sigmoid_prime = 18'b000000010011011000;
		14'b11010101010001:	sigmoid_prime = 18'b000000010011011011;
		14'b11010101010010:	sigmoid_prime = 18'b000000010011011101;
		14'b11010101010011:	sigmoid_prime = 18'b000000010011011111;
		14'b11010101010100:	sigmoid_prime = 18'b000000010011100010;
		14'b11010101010101:	sigmoid_prime = 18'b000000010011100100;
		14'b11010101010110:	sigmoid_prime = 18'b000000010011100111;
		14'b11010101010111:	sigmoid_prime = 18'b000000010011101001;
		14'b11010101011000:	sigmoid_prime = 18'b000000010011101011;
		14'b11010101011001:	sigmoid_prime = 18'b000000010011101110;
		14'b11010101011010:	sigmoid_prime = 18'b000000010011110000;
		14'b11010101011011:	sigmoid_prime = 18'b000000010011110011;
		14'b11010101011100:	sigmoid_prime = 18'b000000010011110101;
		14'b11010101011101:	sigmoid_prime = 18'b000000010011111000;
		14'b11010101011110:	sigmoid_prime = 18'b000000010011111010;
		14'b11010101011111:	sigmoid_prime = 18'b000000010011111101;
		14'b11010101100000:	sigmoid_prime = 18'b000000010011111111;
		14'b11010101100001:	sigmoid_prime = 18'b000000010100000010;
		14'b11010101100010:	sigmoid_prime = 18'b000000010100000100;
		14'b11010101100011:	sigmoid_prime = 18'b000000010100000111;
		14'b11010101100100:	sigmoid_prime = 18'b000000010100001001;
		14'b11010101100101:	sigmoid_prime = 18'b000000010100001100;
		14'b11010101100110:	sigmoid_prime = 18'b000000010100001110;
		14'b11010101100111:	sigmoid_prime = 18'b000000010100010001;
		14'b11010101101000:	sigmoid_prime = 18'b000000010100010011;
		14'b11010101101001:	sigmoid_prime = 18'b000000010100010110;
		14'b11010101101010:	sigmoid_prime = 18'b000000010100011000;
		14'b11010101101011:	sigmoid_prime = 18'b000000010100011011;
		14'b11010101101100:	sigmoid_prime = 18'b000000010100011101;
		14'b11010101101101:	sigmoid_prime = 18'b000000010100100000;
		14'b11010101101110:	sigmoid_prime = 18'b000000010100100010;
		14'b11010101101111:	sigmoid_prime = 18'b000000010100100101;
		14'b11010101110000:	sigmoid_prime = 18'b000000010100100111;
		14'b11010101110001:	sigmoid_prime = 18'b000000010100101010;
		14'b11010101110010:	sigmoid_prime = 18'b000000010100101100;
		14'b11010101110011:	sigmoid_prime = 18'b000000010100101111;
		14'b11010101110100:	sigmoid_prime = 18'b000000010100110010;
		14'b11010101110101:	sigmoid_prime = 18'b000000010100110100;
		14'b11010101110110:	sigmoid_prime = 18'b000000010100110111;
		14'b11010101110111:	sigmoid_prime = 18'b000000010100111001;
		14'b11010101111000:	sigmoid_prime = 18'b000000010100111100;
		14'b11010101111001:	sigmoid_prime = 18'b000000010100111110;
		14'b11010101111010:	sigmoid_prime = 18'b000000010101000001;
		14'b11010101111011:	sigmoid_prime = 18'b000000010101000100;
		14'b11010101111100:	sigmoid_prime = 18'b000000010101000110;
		14'b11010101111101:	sigmoid_prime = 18'b000000010101001001;
		14'b11010101111110:	sigmoid_prime = 18'b000000010101001100;
		14'b11010101111111:	sigmoid_prime = 18'b000000010101001110;
		14'b11010110000000:	sigmoid_prime = 18'b000000010101010001;
		14'b11010110000001:	sigmoid_prime = 18'b000000010101010011;
		14'b11010110000010:	sigmoid_prime = 18'b000000010101010110;
		14'b11010110000011:	sigmoid_prime = 18'b000000010101011001;
		14'b11010110000100:	sigmoid_prime = 18'b000000010101011011;
		14'b11010110000101:	sigmoid_prime = 18'b000000010101011110;
		14'b11010110000110:	sigmoid_prime = 18'b000000010101100001;
		14'b11010110000111:	sigmoid_prime = 18'b000000010101100011;
		14'b11010110001000:	sigmoid_prime = 18'b000000010101100110;
		14'b11010110001001:	sigmoid_prime = 18'b000000010101101001;
		14'b11010110001010:	sigmoid_prime = 18'b000000010101101011;
		14'b11010110001011:	sigmoid_prime = 18'b000000010101101110;
		14'b11010110001100:	sigmoid_prime = 18'b000000010101110001;
		14'b11010110001101:	sigmoid_prime = 18'b000000010101110011;
		14'b11010110001110:	sigmoid_prime = 18'b000000010101110110;
		14'b11010110001111:	sigmoid_prime = 18'b000000010101111001;
		14'b11010110010000:	sigmoid_prime = 18'b000000010101111100;
		14'b11010110010001:	sigmoid_prime = 18'b000000010101111110;
		14'b11010110010010:	sigmoid_prime = 18'b000000010110000001;
		14'b11010110010011:	sigmoid_prime = 18'b000000010110000100;
		14'b11010110010100:	sigmoid_prime = 18'b000000010110000110;
		14'b11010110010101:	sigmoid_prime = 18'b000000010110001001;
		14'b11010110010110:	sigmoid_prime = 18'b000000010110001100;
		14'b11010110010111:	sigmoid_prime = 18'b000000010110001111;
		14'b11010110011000:	sigmoid_prime = 18'b000000010110010001;
		14'b11010110011001:	sigmoid_prime = 18'b000000010110010100;
		14'b11010110011010:	sigmoid_prime = 18'b000000010110010111;
		14'b11010110011011:	sigmoid_prime = 18'b000000010110011010;
		14'b11010110011100:	sigmoid_prime = 18'b000000010110011100;
		14'b11010110011101:	sigmoid_prime = 18'b000000010110011111;
		14'b11010110011110:	sigmoid_prime = 18'b000000010110100010;
		14'b11010110011111:	sigmoid_prime = 18'b000000010110100101;
		14'b11010110100000:	sigmoid_prime = 18'b000000010110101000;
		14'b11010110100001:	sigmoid_prime = 18'b000000010110101010;
		14'b11010110100010:	sigmoid_prime = 18'b000000010110101101;
		14'b11010110100011:	sigmoid_prime = 18'b000000010110110000;
		14'b11010110100100:	sigmoid_prime = 18'b000000010110110011;
		14'b11010110100101:	sigmoid_prime = 18'b000000010110110110;
		14'b11010110100110:	sigmoid_prime = 18'b000000010110111000;
		14'b11010110100111:	sigmoid_prime = 18'b000000010110111011;
		14'b11010110101000:	sigmoid_prime = 18'b000000010110111110;
		14'b11010110101001:	sigmoid_prime = 18'b000000010111000001;
		14'b11010110101010:	sigmoid_prime = 18'b000000010111000100;
		14'b11010110101011:	sigmoid_prime = 18'b000000010111000111;
		14'b11010110101100:	sigmoid_prime = 18'b000000010111001010;
		14'b11010110101101:	sigmoid_prime = 18'b000000010111001100;
		14'b11010110101110:	sigmoid_prime = 18'b000000010111001111;
		14'b11010110101111:	sigmoid_prime = 18'b000000010111010010;
		14'b11010110110000:	sigmoid_prime = 18'b000000010111010101;
		14'b11010110110001:	sigmoid_prime = 18'b000000010111011000;
		14'b11010110110010:	sigmoid_prime = 18'b000000010111011011;
		14'b11010110110011:	sigmoid_prime = 18'b000000010111011110;
		14'b11010110110100:	sigmoid_prime = 18'b000000010111100001;
		14'b11010110110101:	sigmoid_prime = 18'b000000010111100100;
		14'b11010110110110:	sigmoid_prime = 18'b000000010111100110;
		14'b11010110110111:	sigmoid_prime = 18'b000000010111101001;
		14'b11010110111000:	sigmoid_prime = 18'b000000010111101100;
		14'b11010110111001:	sigmoid_prime = 18'b000000010111101111;
		14'b11010110111010:	sigmoid_prime = 18'b000000010111110010;
		14'b11010110111011:	sigmoid_prime = 18'b000000010111110101;
		14'b11010110111100:	sigmoid_prime = 18'b000000010111111000;
		14'b11010110111101:	sigmoid_prime = 18'b000000010111111011;
		14'b11010110111110:	sigmoid_prime = 18'b000000010111111110;
		14'b11010110111111:	sigmoid_prime = 18'b000000011000000001;
		14'b11010111000000:	sigmoid_prime = 18'b000000011000000100;
		14'b11010111000001:	sigmoid_prime = 18'b000000011000000111;
		14'b11010111000010:	sigmoid_prime = 18'b000000011000001010;
		14'b11010111000011:	sigmoid_prime = 18'b000000011000001101;
		14'b11010111000100:	sigmoid_prime = 18'b000000011000010000;
		14'b11010111000101:	sigmoid_prime = 18'b000000011000010011;
		14'b11010111000110:	sigmoid_prime = 18'b000000011000010110;
		14'b11010111000111:	sigmoid_prime = 18'b000000011000011001;
		14'b11010111001000:	sigmoid_prime = 18'b000000011000011100;
		14'b11010111001001:	sigmoid_prime = 18'b000000011000011111;
		14'b11010111001010:	sigmoid_prime = 18'b000000011000100010;
		14'b11010111001011:	sigmoid_prime = 18'b000000011000100101;
		14'b11010111001100:	sigmoid_prime = 18'b000000011000101000;
		14'b11010111001101:	sigmoid_prime = 18'b000000011000101011;
		14'b11010111001110:	sigmoid_prime = 18'b000000011000101110;
		14'b11010111001111:	sigmoid_prime = 18'b000000011000110001;
		14'b11010111010000:	sigmoid_prime = 18'b000000011000110100;
		14'b11010111010001:	sigmoid_prime = 18'b000000011000110111;
		14'b11010111010010:	sigmoid_prime = 18'b000000011000111010;
		14'b11010111010011:	sigmoid_prime = 18'b000000011000111101;
		14'b11010111010100:	sigmoid_prime = 18'b000000011001000000;
		14'b11010111010101:	sigmoid_prime = 18'b000000011001000100;
		14'b11010111010110:	sigmoid_prime = 18'b000000011001000111;
		14'b11010111010111:	sigmoid_prime = 18'b000000011001001010;
		14'b11010111011000:	sigmoid_prime = 18'b000000011001001101;
		14'b11010111011001:	sigmoid_prime = 18'b000000011001010000;
		14'b11010111011010:	sigmoid_prime = 18'b000000011001010011;
		14'b11010111011011:	sigmoid_prime = 18'b000000011001010110;
		14'b11010111011100:	sigmoid_prime = 18'b000000011001011001;
		14'b11010111011101:	sigmoid_prime = 18'b000000011001011101;
		14'b11010111011110:	sigmoid_prime = 18'b000000011001100000;
		14'b11010111011111:	sigmoid_prime = 18'b000000011001100011;
		14'b11010111100000:	sigmoid_prime = 18'b000000011001100110;
		14'b11010111100001:	sigmoid_prime = 18'b000000011001101001;
		14'b11010111100010:	sigmoid_prime = 18'b000000011001101100;
		14'b11010111100011:	sigmoid_prime = 18'b000000011001101111;
		14'b11010111100100:	sigmoid_prime = 18'b000000011001110011;
		14'b11010111100101:	sigmoid_prime = 18'b000000011001110110;
		14'b11010111100110:	sigmoid_prime = 18'b000000011001111001;
		14'b11010111100111:	sigmoid_prime = 18'b000000011001111100;
		14'b11010111101000:	sigmoid_prime = 18'b000000011001111111;
		14'b11010111101001:	sigmoid_prime = 18'b000000011010000011;
		14'b11010111101010:	sigmoid_prime = 18'b000000011010000110;
		14'b11010111101011:	sigmoid_prime = 18'b000000011010001001;
		14'b11010111101100:	sigmoid_prime = 18'b000000011010001100;
		14'b11010111101101:	sigmoid_prime = 18'b000000011010010000;
		14'b11010111101110:	sigmoid_prime = 18'b000000011010010011;
		14'b11010111101111:	sigmoid_prime = 18'b000000011010010110;
		14'b11010111110000:	sigmoid_prime = 18'b000000011010011001;
		14'b11010111110001:	sigmoid_prime = 18'b000000011010011101;
		14'b11010111110010:	sigmoid_prime = 18'b000000011010100000;
		14'b11010111110011:	sigmoid_prime = 18'b000000011010100011;
		14'b11010111110100:	sigmoid_prime = 18'b000000011010100110;
		14'b11010111110101:	sigmoid_prime = 18'b000000011010101010;
		14'b11010111110110:	sigmoid_prime = 18'b000000011010101101;
		14'b11010111110111:	sigmoid_prime = 18'b000000011010110000;
		14'b11010111111000:	sigmoid_prime = 18'b000000011010110100;
		14'b11010111111001:	sigmoid_prime = 18'b000000011010110111;
		14'b11010111111010:	sigmoid_prime = 18'b000000011010111010;
		14'b11010111111011:	sigmoid_prime = 18'b000000011010111110;
		14'b11010111111100:	sigmoid_prime = 18'b000000011011000001;
		14'b11010111111101:	sigmoid_prime = 18'b000000011011000100;
		14'b11010111111110:	sigmoid_prime = 18'b000000011011001000;
		14'b11010111111111:	sigmoid_prime = 18'b000000011011001011;
		14'b11011000000000:	sigmoid_prime = 18'b000000011011001110;
		14'b11011000000001:	sigmoid_prime = 18'b000000011011010010;
		14'b11011000000010:	sigmoid_prime = 18'b000000011011010101;
		14'b11011000000011:	sigmoid_prime = 18'b000000011011011000;
		14'b11011000000100:	sigmoid_prime = 18'b000000011011011100;
		14'b11011000000101:	sigmoid_prime = 18'b000000011011011111;
		14'b11011000000110:	sigmoid_prime = 18'b000000011011100011;
		14'b11011000000111:	sigmoid_prime = 18'b000000011011100110;
		14'b11011000001000:	sigmoid_prime = 18'b000000011011101001;
		14'b11011000001001:	sigmoid_prime = 18'b000000011011101101;
		14'b11011000001010:	sigmoid_prime = 18'b000000011011110000;
		14'b11011000001011:	sigmoid_prime = 18'b000000011011110100;
		14'b11011000001100:	sigmoid_prime = 18'b000000011011110111;
		14'b11011000001101:	sigmoid_prime = 18'b000000011011111010;
		14'b11011000001110:	sigmoid_prime = 18'b000000011011111110;
		14'b11011000001111:	sigmoid_prime = 18'b000000011100000001;
		14'b11011000010000:	sigmoid_prime = 18'b000000011100000101;
		14'b11011000010001:	sigmoid_prime = 18'b000000011100001000;
		14'b11011000010010:	sigmoid_prime = 18'b000000011100001100;
		14'b11011000010011:	sigmoid_prime = 18'b000000011100001111;
		14'b11011000010100:	sigmoid_prime = 18'b000000011100010011;
		14'b11011000010101:	sigmoid_prime = 18'b000000011100010110;
		14'b11011000010110:	sigmoid_prime = 18'b000000011100011010;
		14'b11011000010111:	sigmoid_prime = 18'b000000011100011101;
		14'b11011000011000:	sigmoid_prime = 18'b000000011100100001;
		14'b11011000011001:	sigmoid_prime = 18'b000000011100100100;
		14'b11011000011010:	sigmoid_prime = 18'b000000011100101000;
		14'b11011000011011:	sigmoid_prime = 18'b000000011100101011;
		14'b11011000011100:	sigmoid_prime = 18'b000000011100101111;
		14'b11011000011101:	sigmoid_prime = 18'b000000011100110010;
		14'b11011000011110:	sigmoid_prime = 18'b000000011100110110;
		14'b11011000011111:	sigmoid_prime = 18'b000000011100111001;
		14'b11011000100000:	sigmoid_prime = 18'b000000011100111101;
		14'b11011000100001:	sigmoid_prime = 18'b000000011101000001;
		14'b11011000100010:	sigmoid_prime = 18'b000000011101000100;
		14'b11011000100011:	sigmoid_prime = 18'b000000011101001000;
		14'b11011000100100:	sigmoid_prime = 18'b000000011101001011;
		14'b11011000100101:	sigmoid_prime = 18'b000000011101001111;
		14'b11011000100110:	sigmoid_prime = 18'b000000011101010011;
		14'b11011000100111:	sigmoid_prime = 18'b000000011101010110;
		14'b11011000101000:	sigmoid_prime = 18'b000000011101011010;
		14'b11011000101001:	sigmoid_prime = 18'b000000011101011101;
		14'b11011000101010:	sigmoid_prime = 18'b000000011101100001;
		14'b11011000101011:	sigmoid_prime = 18'b000000011101100101;
		14'b11011000101100:	sigmoid_prime = 18'b000000011101101000;
		14'b11011000101101:	sigmoid_prime = 18'b000000011101101100;
		14'b11011000101110:	sigmoid_prime = 18'b000000011101110000;
		14'b11011000101111:	sigmoid_prime = 18'b000000011101110011;
		14'b11011000110000:	sigmoid_prime = 18'b000000011101110111;
		14'b11011000110001:	sigmoid_prime = 18'b000000011101111011;
		14'b11011000110010:	sigmoid_prime = 18'b000000011101111110;
		14'b11011000110011:	sigmoid_prime = 18'b000000011110000010;
		14'b11011000110100:	sigmoid_prime = 18'b000000011110000110;
		14'b11011000110101:	sigmoid_prime = 18'b000000011110001001;
		14'b11011000110110:	sigmoid_prime = 18'b000000011110001101;
		14'b11011000110111:	sigmoid_prime = 18'b000000011110010001;
		14'b11011000111000:	sigmoid_prime = 18'b000000011110010101;
		14'b11011000111001:	sigmoid_prime = 18'b000000011110011000;
		14'b11011000111010:	sigmoid_prime = 18'b000000011110011100;
		14'b11011000111011:	sigmoid_prime = 18'b000000011110100000;
		14'b11011000111100:	sigmoid_prime = 18'b000000011110100100;
		14'b11011000111101:	sigmoid_prime = 18'b000000011110100111;
		14'b11011000111110:	sigmoid_prime = 18'b000000011110101011;
		14'b11011000111111:	sigmoid_prime = 18'b000000011110101111;
		14'b11011001000000:	sigmoid_prime = 18'b000000011110110011;
		14'b11011001000001:	sigmoid_prime = 18'b000000011110110111;
		14'b11011001000010:	sigmoid_prime = 18'b000000011110111010;
		14'b11011001000011:	sigmoid_prime = 18'b000000011110111110;
		14'b11011001000100:	sigmoid_prime = 18'b000000011111000010;
		14'b11011001000101:	sigmoid_prime = 18'b000000011111000110;
		14'b11011001000110:	sigmoid_prime = 18'b000000011111001010;
		14'b11011001000111:	sigmoid_prime = 18'b000000011111001101;
		14'b11011001001000:	sigmoid_prime = 18'b000000011111010001;
		14'b11011001001001:	sigmoid_prime = 18'b000000011111010101;
		14'b11011001001010:	sigmoid_prime = 18'b000000011111011001;
		14'b11011001001011:	sigmoid_prime = 18'b000000011111011101;
		14'b11011001001100:	sigmoid_prime = 18'b000000011111100001;
		14'b11011001001101:	sigmoid_prime = 18'b000000011111100101;
		14'b11011001001110:	sigmoid_prime = 18'b000000011111101001;
		14'b11011001001111:	sigmoid_prime = 18'b000000011111101100;
		14'b11011001010000:	sigmoid_prime = 18'b000000011111110000;
		14'b11011001010001:	sigmoid_prime = 18'b000000011111110100;
		14'b11011001010010:	sigmoid_prime = 18'b000000011111111000;
		14'b11011001010011:	sigmoid_prime = 18'b000000011111111100;
		14'b11011001010100:	sigmoid_prime = 18'b000000100000000000;
		14'b11011001010101:	sigmoid_prime = 18'b000000100000000100;
		14'b11011001010110:	sigmoid_prime = 18'b000000100000001000;
		14'b11011001010111:	sigmoid_prime = 18'b000000100000001100;
		14'b11011001011000:	sigmoid_prime = 18'b000000100000010000;
		14'b11011001011001:	sigmoid_prime = 18'b000000100000010100;
		14'b11011001011010:	sigmoid_prime = 18'b000000100000011000;
		14'b11011001011011:	sigmoid_prime = 18'b000000100000011100;
		14'b11011001011100:	sigmoid_prime = 18'b000000100000100000;
		14'b11011001011101:	sigmoid_prime = 18'b000000100000100100;
		14'b11011001011110:	sigmoid_prime = 18'b000000100000101000;
		14'b11011001011111:	sigmoid_prime = 18'b000000100000101100;
		14'b11011001100000:	sigmoid_prime = 18'b000000100000110000;
		14'b11011001100001:	sigmoid_prime = 18'b000000100000110100;
		14'b11011001100010:	sigmoid_prime = 18'b000000100000111000;
		14'b11011001100011:	sigmoid_prime = 18'b000000100000111100;
		14'b11011001100100:	sigmoid_prime = 18'b000000100001000000;
		14'b11011001100101:	sigmoid_prime = 18'b000000100001000100;
		14'b11011001100110:	sigmoid_prime = 18'b000000100001001000;
		14'b11011001100111:	sigmoid_prime = 18'b000000100001001100;
		14'b11011001101000:	sigmoid_prime = 18'b000000100001010000;
		14'b11011001101001:	sigmoid_prime = 18'b000000100001010100;
		14'b11011001101010:	sigmoid_prime = 18'b000000100001011001;
		14'b11011001101011:	sigmoid_prime = 18'b000000100001011101;
		14'b11011001101100:	sigmoid_prime = 18'b000000100001100001;
		14'b11011001101101:	sigmoid_prime = 18'b000000100001100101;
		14'b11011001101110:	sigmoid_prime = 18'b000000100001101001;
		14'b11011001101111:	sigmoid_prime = 18'b000000100001101101;
		14'b11011001110000:	sigmoid_prime = 18'b000000100001110001;
		14'b11011001110001:	sigmoid_prime = 18'b000000100001110101;
		14'b11011001110010:	sigmoid_prime = 18'b000000100001111010;
		14'b11011001110011:	sigmoid_prime = 18'b000000100001111110;
		14'b11011001110100:	sigmoid_prime = 18'b000000100010000010;
		14'b11011001110101:	sigmoid_prime = 18'b000000100010000110;
		14'b11011001110110:	sigmoid_prime = 18'b000000100010001010;
		14'b11011001110111:	sigmoid_prime = 18'b000000100010001111;
		14'b11011001111000:	sigmoid_prime = 18'b000000100010010011;
		14'b11011001111001:	sigmoid_prime = 18'b000000100010010111;
		14'b11011001111010:	sigmoid_prime = 18'b000000100010011011;
		14'b11011001111011:	sigmoid_prime = 18'b000000100010011111;
		14'b11011001111100:	sigmoid_prime = 18'b000000100010100100;
		14'b11011001111101:	sigmoid_prime = 18'b000000100010101000;
		14'b11011001111110:	sigmoid_prime = 18'b000000100010101100;
		14'b11011001111111:	sigmoid_prime = 18'b000000100010110000;
		14'b11011010000000:	sigmoid_prime = 18'b000000100010110101;
		14'b11011010000001:	sigmoid_prime = 18'b000000100010111001;
		14'b11011010000010:	sigmoid_prime = 18'b000000100010111101;
		14'b11011010000011:	sigmoid_prime = 18'b000000100011000010;
		14'b11011010000100:	sigmoid_prime = 18'b000000100011000110;
		14'b11011010000101:	sigmoid_prime = 18'b000000100011001010;
		14'b11011010000110:	sigmoid_prime = 18'b000000100011001111;
		14'b11011010000111:	sigmoid_prime = 18'b000000100011010011;
		14'b11011010001000:	sigmoid_prime = 18'b000000100011010111;
		14'b11011010001001:	sigmoid_prime = 18'b000000100011011100;
		14'b11011010001010:	sigmoid_prime = 18'b000000100011100000;
		14'b11011010001011:	sigmoid_prime = 18'b000000100011100100;
		14'b11011010001100:	sigmoid_prime = 18'b000000100011101001;
		14'b11011010001101:	sigmoid_prime = 18'b000000100011101101;
		14'b11011010001110:	sigmoid_prime = 18'b000000100011110001;
		14'b11011010001111:	sigmoid_prime = 18'b000000100011110110;
		14'b11011010010000:	sigmoid_prime = 18'b000000100011111010;
		14'b11011010010001:	sigmoid_prime = 18'b000000100011111111;
		14'b11011010010010:	sigmoid_prime = 18'b000000100100000011;
		14'b11011010010011:	sigmoid_prime = 18'b000000100100001000;
		14'b11011010010100:	sigmoid_prime = 18'b000000100100001100;
		14'b11011010010101:	sigmoid_prime = 18'b000000100100010000;
		14'b11011010010110:	sigmoid_prime = 18'b000000100100010101;
		14'b11011010010111:	sigmoid_prime = 18'b000000100100011001;
		14'b11011010011000:	sigmoid_prime = 18'b000000100100011110;
		14'b11011010011001:	sigmoid_prime = 18'b000000100100100010;
		14'b11011010011010:	sigmoid_prime = 18'b000000100100100111;
		14'b11011010011011:	sigmoid_prime = 18'b000000100100101011;
		14'b11011010011100:	sigmoid_prime = 18'b000000100100110000;
		14'b11011010011101:	sigmoid_prime = 18'b000000100100110100;
		14'b11011010011110:	sigmoid_prime = 18'b000000100100111001;
		14'b11011010011111:	sigmoid_prime = 18'b000000100100111101;
		14'b11011010100000:	sigmoid_prime = 18'b000000100101000010;
		14'b11011010100001:	sigmoid_prime = 18'b000000100101000110;
		14'b11011010100010:	sigmoid_prime = 18'b000000100101001011;
		14'b11011010100011:	sigmoid_prime = 18'b000000100101010000;
		14'b11011010100100:	sigmoid_prime = 18'b000000100101010100;
		14'b11011010100101:	sigmoid_prime = 18'b000000100101011001;
		14'b11011010100110:	sigmoid_prime = 18'b000000100101011101;
		14'b11011010100111:	sigmoid_prime = 18'b000000100101100010;
		14'b11011010101000:	sigmoid_prime = 18'b000000100101100111;
		14'b11011010101001:	sigmoid_prime = 18'b000000100101101011;
		14'b11011010101010:	sigmoid_prime = 18'b000000100101110000;
		14'b11011010101011:	sigmoid_prime = 18'b000000100101110100;
		14'b11011010101100:	sigmoid_prime = 18'b000000100101111001;
		14'b11011010101101:	sigmoid_prime = 18'b000000100101111110;
		14'b11011010101110:	sigmoid_prime = 18'b000000100110000010;
		14'b11011010101111:	sigmoid_prime = 18'b000000100110000111;
		14'b11011010110000:	sigmoid_prime = 18'b000000100110001100;
		14'b11011010110001:	sigmoid_prime = 18'b000000100110010000;
		14'b11011010110010:	sigmoid_prime = 18'b000000100110010101;
		14'b11011010110011:	sigmoid_prime = 18'b000000100110011010;
		14'b11011010110100:	sigmoid_prime = 18'b000000100110011111;
		14'b11011010110101:	sigmoid_prime = 18'b000000100110100011;
		14'b11011010110110:	sigmoid_prime = 18'b000000100110101000;
		14'b11011010110111:	sigmoid_prime = 18'b000000100110101101;
		14'b11011010111000:	sigmoid_prime = 18'b000000100110110001;
		14'b11011010111001:	sigmoid_prime = 18'b000000100110110110;
		14'b11011010111010:	sigmoid_prime = 18'b000000100110111011;
		14'b11011010111011:	sigmoid_prime = 18'b000000100111000000;
		14'b11011010111100:	sigmoid_prime = 18'b000000100111000101;
		14'b11011010111101:	sigmoid_prime = 18'b000000100111001001;
		14'b11011010111110:	sigmoid_prime = 18'b000000100111001110;
		14'b11011010111111:	sigmoid_prime = 18'b000000100111010011;
		14'b11011011000000:	sigmoid_prime = 18'b000000100111011000;
		14'b11011011000001:	sigmoid_prime = 18'b000000100111011101;
		14'b11011011000010:	sigmoid_prime = 18'b000000100111100001;
		14'b11011011000011:	sigmoid_prime = 18'b000000100111100110;
		14'b11011011000100:	sigmoid_prime = 18'b000000100111101011;
		14'b11011011000101:	sigmoid_prime = 18'b000000100111110000;
		14'b11011011000110:	sigmoid_prime = 18'b000000100111110101;
		14'b11011011000111:	sigmoid_prime = 18'b000000100111111010;
		14'b11011011001000:	sigmoid_prime = 18'b000000100111111111;
		14'b11011011001001:	sigmoid_prime = 18'b000000101000000100;
		14'b11011011001010:	sigmoid_prime = 18'b000000101000001001;
		14'b11011011001011:	sigmoid_prime = 18'b000000101000001101;
		14'b11011011001100:	sigmoid_prime = 18'b000000101000010010;
		14'b11011011001101:	sigmoid_prime = 18'b000000101000010111;
		14'b11011011001110:	sigmoid_prime = 18'b000000101000011100;
		14'b11011011001111:	sigmoid_prime = 18'b000000101000100001;
		14'b11011011010000:	sigmoid_prime = 18'b000000101000100110;
		14'b11011011010001:	sigmoid_prime = 18'b000000101000101011;
		14'b11011011010010:	sigmoid_prime = 18'b000000101000110000;
		14'b11011011010011:	sigmoid_prime = 18'b000000101000110101;
		14'b11011011010100:	sigmoid_prime = 18'b000000101000111010;
		14'b11011011010101:	sigmoid_prime = 18'b000000101000111111;
		14'b11011011010110:	sigmoid_prime = 18'b000000101001000100;
		14'b11011011010111:	sigmoid_prime = 18'b000000101001001001;
		14'b11011011011000:	sigmoid_prime = 18'b000000101001001110;
		14'b11011011011001:	sigmoid_prime = 18'b000000101001010011;
		14'b11011011011010:	sigmoid_prime = 18'b000000101001011000;
		14'b11011011011011:	sigmoid_prime = 18'b000000101001011101;
		14'b11011011011100:	sigmoid_prime = 18'b000000101001100011;
		14'b11011011011101:	sigmoid_prime = 18'b000000101001101000;
		14'b11011011011110:	sigmoid_prime = 18'b000000101001101101;
		14'b11011011011111:	sigmoid_prime = 18'b000000101001110010;
		14'b11011011100000:	sigmoid_prime = 18'b000000101001110111;
		14'b11011011100001:	sigmoid_prime = 18'b000000101001111100;
		14'b11011011100010:	sigmoid_prime = 18'b000000101010000001;
		14'b11011011100011:	sigmoid_prime = 18'b000000101010000110;
		14'b11011011100100:	sigmoid_prime = 18'b000000101010001100;
		14'b11011011100101:	sigmoid_prime = 18'b000000101010010001;
		14'b11011011100110:	sigmoid_prime = 18'b000000101010010110;
		14'b11011011100111:	sigmoid_prime = 18'b000000101010011011;
		14'b11011011101000:	sigmoid_prime = 18'b000000101010100000;
		14'b11011011101001:	sigmoid_prime = 18'b000000101010100110;
		14'b11011011101010:	sigmoid_prime = 18'b000000101010101011;
		14'b11011011101011:	sigmoid_prime = 18'b000000101010110000;
		14'b11011011101100:	sigmoid_prime = 18'b000000101010110101;
		14'b11011011101101:	sigmoid_prime = 18'b000000101010111010;
		14'b11011011101110:	sigmoid_prime = 18'b000000101011000000;
		14'b11011011101111:	sigmoid_prime = 18'b000000101011000101;
		14'b11011011110000:	sigmoid_prime = 18'b000000101011001010;
		14'b11011011110001:	sigmoid_prime = 18'b000000101011010000;
		14'b11011011110010:	sigmoid_prime = 18'b000000101011010101;
		14'b11011011110011:	sigmoid_prime = 18'b000000101011011010;
		14'b11011011110100:	sigmoid_prime = 18'b000000101011011111;
		14'b11011011110101:	sigmoid_prime = 18'b000000101011100101;
		14'b11011011110110:	sigmoid_prime = 18'b000000101011101010;
		14'b11011011110111:	sigmoid_prime = 18'b000000101011101111;
		14'b11011011111000:	sigmoid_prime = 18'b000000101011110101;
		14'b11011011111001:	sigmoid_prime = 18'b000000101011111010;
		14'b11011011111010:	sigmoid_prime = 18'b000000101100000000;
		14'b11011011111011:	sigmoid_prime = 18'b000000101100000101;
		14'b11011011111100:	sigmoid_prime = 18'b000000101100001010;
		14'b11011011111101:	sigmoid_prime = 18'b000000101100010000;
		14'b11011011111110:	sigmoid_prime = 18'b000000101100010101;
		14'b11011011111111:	sigmoid_prime = 18'b000000101100011011;
		14'b11011100000000:	sigmoid_prime = 18'b000000101100100000;
		14'b11011100000001:	sigmoid_prime = 18'b000000101100100101;
		14'b11011100000010:	sigmoid_prime = 18'b000000101100101011;
		14'b11011100000011:	sigmoid_prime = 18'b000000101100110000;
		14'b11011100000100:	sigmoid_prime = 18'b000000101100110110;
		14'b11011100000101:	sigmoid_prime = 18'b000000101100111011;
		14'b11011100000110:	sigmoid_prime = 18'b000000101101000001;
		14'b11011100000111:	sigmoid_prime = 18'b000000101101000110;
		14'b11011100001000:	sigmoid_prime = 18'b000000101101001100;
		14'b11011100001001:	sigmoid_prime = 18'b000000101101010001;
		14'b11011100001010:	sigmoid_prime = 18'b000000101101010111;
		14'b11011100001011:	sigmoid_prime = 18'b000000101101011100;
		14'b11011100001100:	sigmoid_prime = 18'b000000101101100010;
		14'b11011100001101:	sigmoid_prime = 18'b000000101101101000;
		14'b11011100001110:	sigmoid_prime = 18'b000000101101101101;
		14'b11011100001111:	sigmoid_prime = 18'b000000101101110011;
		14'b11011100010000:	sigmoid_prime = 18'b000000101101111000;
		14'b11011100010001:	sigmoid_prime = 18'b000000101101111110;
		14'b11011100010010:	sigmoid_prime = 18'b000000101110000100;
		14'b11011100010011:	sigmoid_prime = 18'b000000101110001001;
		14'b11011100010100:	sigmoid_prime = 18'b000000101110001111;
		14'b11011100010101:	sigmoid_prime = 18'b000000101110010101;
		14'b11011100010110:	sigmoid_prime = 18'b000000101110011010;
		14'b11011100010111:	sigmoid_prime = 18'b000000101110100000;
		14'b11011100011000:	sigmoid_prime = 18'b000000101110100110;
		14'b11011100011001:	sigmoid_prime = 18'b000000101110101011;
		14'b11011100011010:	sigmoid_prime = 18'b000000101110110001;
		14'b11011100011011:	sigmoid_prime = 18'b000000101110110111;
		14'b11011100011100:	sigmoid_prime = 18'b000000101110111100;
		14'b11011100011101:	sigmoid_prime = 18'b000000101111000010;
		14'b11011100011110:	sigmoid_prime = 18'b000000101111001000;
		14'b11011100011111:	sigmoid_prime = 18'b000000101111001110;
		14'b11011100100000:	sigmoid_prime = 18'b000000101111010011;
		14'b11011100100001:	sigmoid_prime = 18'b000000101111011001;
		14'b11011100100010:	sigmoid_prime = 18'b000000101111011111;
		14'b11011100100011:	sigmoid_prime = 18'b000000101111100101;
		14'b11011100100100:	sigmoid_prime = 18'b000000101111101011;
		14'b11011100100101:	sigmoid_prime = 18'b000000101111110000;
		14'b11011100100110:	sigmoid_prime = 18'b000000101111110110;
		14'b11011100100111:	sigmoid_prime = 18'b000000101111111100;
		14'b11011100101000:	sigmoid_prime = 18'b000000110000000010;
		14'b11011100101001:	sigmoid_prime = 18'b000000110000001000;
		14'b11011100101010:	sigmoid_prime = 18'b000000110000001110;
		14'b11011100101011:	sigmoid_prime = 18'b000000110000010100;
		14'b11011100101100:	sigmoid_prime = 18'b000000110000011010;
		14'b11011100101101:	sigmoid_prime = 18'b000000110000011111;
		14'b11011100101110:	sigmoid_prime = 18'b000000110000100101;
		14'b11011100101111:	sigmoid_prime = 18'b000000110000101011;
		14'b11011100110000:	sigmoid_prime = 18'b000000110000110001;
		14'b11011100110001:	sigmoid_prime = 18'b000000110000110111;
		14'b11011100110010:	sigmoid_prime = 18'b000000110000111101;
		14'b11011100110011:	sigmoid_prime = 18'b000000110001000011;
		14'b11011100110100:	sigmoid_prime = 18'b000000110001001001;
		14'b11011100110101:	sigmoid_prime = 18'b000000110001001111;
		14'b11011100110110:	sigmoid_prime = 18'b000000110001010101;
		14'b11011100110111:	sigmoid_prime = 18'b000000110001011011;
		14'b11011100111000:	sigmoid_prime = 18'b000000110001100001;
		14'b11011100111001:	sigmoid_prime = 18'b000000110001100111;
		14'b11011100111010:	sigmoid_prime = 18'b000000110001101101;
		14'b11011100111011:	sigmoid_prime = 18'b000000110001110011;
		14'b11011100111100:	sigmoid_prime = 18'b000000110001111001;
		14'b11011100111101:	sigmoid_prime = 18'b000000110010000000;
		14'b11011100111110:	sigmoid_prime = 18'b000000110010000110;
		14'b11011100111111:	sigmoid_prime = 18'b000000110010001100;
		14'b11011101000000:	sigmoid_prime = 18'b000000110010010010;
		14'b11011101000001:	sigmoid_prime = 18'b000000110010011000;
		14'b11011101000010:	sigmoid_prime = 18'b000000110010011110;
		14'b11011101000011:	sigmoid_prime = 18'b000000110010100100;
		14'b11011101000100:	sigmoid_prime = 18'b000000110010101010;
		14'b11011101000101:	sigmoid_prime = 18'b000000110010110001;
		14'b11011101000110:	sigmoid_prime = 18'b000000110010110111;
		14'b11011101000111:	sigmoid_prime = 18'b000000110010111101;
		14'b11011101001000:	sigmoid_prime = 18'b000000110011000011;
		14'b11011101001001:	sigmoid_prime = 18'b000000110011001001;
		14'b11011101001010:	sigmoid_prime = 18'b000000110011010000;
		14'b11011101001011:	sigmoid_prime = 18'b000000110011010110;
		14'b11011101001100:	sigmoid_prime = 18'b000000110011011100;
		14'b11011101001101:	sigmoid_prime = 18'b000000110011100011;
		14'b11011101001110:	sigmoid_prime = 18'b000000110011101001;
		14'b11011101001111:	sigmoid_prime = 18'b000000110011101111;
		14'b11011101010000:	sigmoid_prime = 18'b000000110011110101;
		14'b11011101010001:	sigmoid_prime = 18'b000000110011111100;
		14'b11011101010010:	sigmoid_prime = 18'b000000110100000010;
		14'b11011101010011:	sigmoid_prime = 18'b000000110100001000;
		14'b11011101010100:	sigmoid_prime = 18'b000000110100001111;
		14'b11011101010101:	sigmoid_prime = 18'b000000110100010101;
		14'b11011101010110:	sigmoid_prime = 18'b000000110100011100;
		14'b11011101010111:	sigmoid_prime = 18'b000000110100100010;
		14'b11011101011000:	sigmoid_prime = 18'b000000110100101000;
		14'b11011101011001:	sigmoid_prime = 18'b000000110100101111;
		14'b11011101011010:	sigmoid_prime = 18'b000000110100110101;
		14'b11011101011011:	sigmoid_prime = 18'b000000110100111100;
		14'b11011101011100:	sigmoid_prime = 18'b000000110101000010;
		14'b11011101011101:	sigmoid_prime = 18'b000000110101001000;
		14'b11011101011110:	sigmoid_prime = 18'b000000110101001111;
		14'b11011101011111:	sigmoid_prime = 18'b000000110101010101;
		14'b11011101100000:	sigmoid_prime = 18'b000000110101011100;
		14'b11011101100001:	sigmoid_prime = 18'b000000110101100010;
		14'b11011101100010:	sigmoid_prime = 18'b000000110101101001;
		14'b11011101100011:	sigmoid_prime = 18'b000000110101110000;
		14'b11011101100100:	sigmoid_prime = 18'b000000110101110110;
		14'b11011101100101:	sigmoid_prime = 18'b000000110101111101;
		14'b11011101100110:	sigmoid_prime = 18'b000000110110000011;
		14'b11011101100111:	sigmoid_prime = 18'b000000110110001010;
		14'b11011101101000:	sigmoid_prime = 18'b000000110110010000;
		14'b11011101101001:	sigmoid_prime = 18'b000000110110010111;
		14'b11011101101010:	sigmoid_prime = 18'b000000110110011110;
		14'b11011101101011:	sigmoid_prime = 18'b000000110110100100;
		14'b11011101101100:	sigmoid_prime = 18'b000000110110101011;
		14'b11011101101101:	sigmoid_prime = 18'b000000110110110010;
		14'b11011101101110:	sigmoid_prime = 18'b000000110110111000;
		14'b11011101101111:	sigmoid_prime = 18'b000000110110111111;
		14'b11011101110000:	sigmoid_prime = 18'b000000110111000110;
		14'b11011101110001:	sigmoid_prime = 18'b000000110111001100;
		14'b11011101110010:	sigmoid_prime = 18'b000000110111010011;
		14'b11011101110011:	sigmoid_prime = 18'b000000110111011010;
		14'b11011101110100:	sigmoid_prime = 18'b000000110111100000;
		14'b11011101110101:	sigmoid_prime = 18'b000000110111100111;
		14'b11011101110110:	sigmoid_prime = 18'b000000110111101110;
		14'b11011101110111:	sigmoid_prime = 18'b000000110111110101;
		14'b11011101111000:	sigmoid_prime = 18'b000000110111111100;
		14'b11011101111001:	sigmoid_prime = 18'b000000111000000010;
		14'b11011101111010:	sigmoid_prime = 18'b000000111000001001;
		14'b11011101111011:	sigmoid_prime = 18'b000000111000010000;
		14'b11011101111100:	sigmoid_prime = 18'b000000111000010111;
		14'b11011101111101:	sigmoid_prime = 18'b000000111000011110;
		14'b11011101111110:	sigmoid_prime = 18'b000000111000100101;
		14'b11011101111111:	sigmoid_prime = 18'b000000111000101011;
		14'b11011110000000:	sigmoid_prime = 18'b000000111000110010;
		14'b11011110000001:	sigmoid_prime = 18'b000000111000111001;
		14'b11011110000010:	sigmoid_prime = 18'b000000111001000000;
		14'b11011110000011:	sigmoid_prime = 18'b000000111001000111;
		14'b11011110000100:	sigmoid_prime = 18'b000000111001001110;
		14'b11011110000101:	sigmoid_prime = 18'b000000111001010101;
		14'b11011110000110:	sigmoid_prime = 18'b000000111001011100;
		14'b11011110000111:	sigmoid_prime = 18'b000000111001100011;
		14'b11011110001000:	sigmoid_prime = 18'b000000111001101010;
		14'b11011110001001:	sigmoid_prime = 18'b000000111001110001;
		14'b11011110001010:	sigmoid_prime = 18'b000000111001111000;
		14'b11011110001011:	sigmoid_prime = 18'b000000111001111111;
		14'b11011110001100:	sigmoid_prime = 18'b000000111010000110;
		14'b11011110001101:	sigmoid_prime = 18'b000000111010001101;
		14'b11011110001110:	sigmoid_prime = 18'b000000111010010100;
		14'b11011110001111:	sigmoid_prime = 18'b000000111010011011;
		14'b11011110010000:	sigmoid_prime = 18'b000000111010100010;
		14'b11011110010001:	sigmoid_prime = 18'b000000111010101001;
		14'b11011110010010:	sigmoid_prime = 18'b000000111010110001;
		14'b11011110010011:	sigmoid_prime = 18'b000000111010111000;
		14'b11011110010100:	sigmoid_prime = 18'b000000111010111111;
		14'b11011110010101:	sigmoid_prime = 18'b000000111011000110;
		14'b11011110010110:	sigmoid_prime = 18'b000000111011001101;
		14'b11011110010111:	sigmoid_prime = 18'b000000111011010100;
		14'b11011110011000:	sigmoid_prime = 18'b000000111011011100;
		14'b11011110011001:	sigmoid_prime = 18'b000000111011100011;
		14'b11011110011010:	sigmoid_prime = 18'b000000111011101010;
		14'b11011110011011:	sigmoid_prime = 18'b000000111011110001;
		14'b11011110011100:	sigmoid_prime = 18'b000000111011111001;
		14'b11011110011101:	sigmoid_prime = 18'b000000111100000000;
		14'b11011110011110:	sigmoid_prime = 18'b000000111100000111;
		14'b11011110011111:	sigmoid_prime = 18'b000000111100001110;
		14'b11011110100000:	sigmoid_prime = 18'b000000111100010110;
		14'b11011110100001:	sigmoid_prime = 18'b000000111100011101;
		14'b11011110100010:	sigmoid_prime = 18'b000000111100100100;
		14'b11011110100011:	sigmoid_prime = 18'b000000111100101100;
		14'b11011110100100:	sigmoid_prime = 18'b000000111100110011;
		14'b11011110100101:	sigmoid_prime = 18'b000000111100111011;
		14'b11011110100110:	sigmoid_prime = 18'b000000111101000010;
		14'b11011110100111:	sigmoid_prime = 18'b000000111101001001;
		14'b11011110101000:	sigmoid_prime = 18'b000000111101010001;
		14'b11011110101001:	sigmoid_prime = 18'b000000111101011000;
		14'b11011110101010:	sigmoid_prime = 18'b000000111101100000;
		14'b11011110101011:	sigmoid_prime = 18'b000000111101100111;
		14'b11011110101100:	sigmoid_prime = 18'b000000111101101111;
		14'b11011110101101:	sigmoid_prime = 18'b000000111101110110;
		14'b11011110101110:	sigmoid_prime = 18'b000000111101111110;
		14'b11011110101111:	sigmoid_prime = 18'b000000111110000101;
		14'b11011110110000:	sigmoid_prime = 18'b000000111110001101;
		14'b11011110110001:	sigmoid_prime = 18'b000000111110010100;
		14'b11011110110010:	sigmoid_prime = 18'b000000111110011100;
		14'b11011110110011:	sigmoid_prime = 18'b000000111110100011;
		14'b11011110110100:	sigmoid_prime = 18'b000000111110101011;
		14'b11011110110101:	sigmoid_prime = 18'b000000111110110010;
		14'b11011110110110:	sigmoid_prime = 18'b000000111110111010;
		14'b11011110110111:	sigmoid_prime = 18'b000000111111000010;
		14'b11011110111000:	sigmoid_prime = 18'b000000111111001001;
		14'b11011110111001:	sigmoid_prime = 18'b000000111111010001;
		14'b11011110111010:	sigmoid_prime = 18'b000000111111011001;
		14'b11011110111011:	sigmoid_prime = 18'b000000111111100000;
		14'b11011110111100:	sigmoid_prime = 18'b000000111111101000;
		14'b11011110111101:	sigmoid_prime = 18'b000000111111110000;
		14'b11011110111110:	sigmoid_prime = 18'b000000111111110111;
		14'b11011110111111:	sigmoid_prime = 18'b000000111111111111;
		14'b11011111000000:	sigmoid_prime = 18'b000001000000000111;
		14'b11011111000001:	sigmoid_prime = 18'b000001000000001111;
		14'b11011111000010:	sigmoid_prime = 18'b000001000000010110;
		14'b11011111000011:	sigmoid_prime = 18'b000001000000011110;
		14'b11011111000100:	sigmoid_prime = 18'b000001000000100110;
		14'b11011111000101:	sigmoid_prime = 18'b000001000000101110;
		14'b11011111000110:	sigmoid_prime = 18'b000001000000110110;
		14'b11011111000111:	sigmoid_prime = 18'b000001000000111110;
		14'b11011111001000:	sigmoid_prime = 18'b000001000001000101;
		14'b11011111001001:	sigmoid_prime = 18'b000001000001001101;
		14'b11011111001010:	sigmoid_prime = 18'b000001000001010101;
		14'b11011111001011:	sigmoid_prime = 18'b000001000001011101;
		14'b11011111001100:	sigmoid_prime = 18'b000001000001100101;
		14'b11011111001101:	sigmoid_prime = 18'b000001000001101101;
		14'b11011111001110:	sigmoid_prime = 18'b000001000001110101;
		14'b11011111001111:	sigmoid_prime = 18'b000001000001111101;
		14'b11011111010000:	sigmoid_prime = 18'b000001000010000101;
		14'b11011111010001:	sigmoid_prime = 18'b000001000010001101;
		14'b11011111010010:	sigmoid_prime = 18'b000001000010010101;
		14'b11011111010011:	sigmoid_prime = 18'b000001000010011101;
		14'b11011111010100:	sigmoid_prime = 18'b000001000010100101;
		14'b11011111010101:	sigmoid_prime = 18'b000001000010101101;
		14'b11011111010110:	sigmoid_prime = 18'b000001000010110101;
		14'b11011111010111:	sigmoid_prime = 18'b000001000010111101;
		14'b11011111011000:	sigmoid_prime = 18'b000001000011000101;
		14'b11011111011001:	sigmoid_prime = 18'b000001000011001101;
		14'b11011111011010:	sigmoid_prime = 18'b000001000011010110;
		14'b11011111011011:	sigmoid_prime = 18'b000001000011011110;
		14'b11011111011100:	sigmoid_prime = 18'b000001000011100110;
		14'b11011111011101:	sigmoid_prime = 18'b000001000011101110;
		14'b11011111011110:	sigmoid_prime = 18'b000001000011110110;
		14'b11011111011111:	sigmoid_prime = 18'b000001000011111110;
		14'b11011111100000:	sigmoid_prime = 18'b000001000100000111;
		14'b11011111100001:	sigmoid_prime = 18'b000001000100001111;
		14'b11011111100010:	sigmoid_prime = 18'b000001000100010111;
		14'b11011111100011:	sigmoid_prime = 18'b000001000100011111;
		14'b11011111100100:	sigmoid_prime = 18'b000001000100101000;
		14'b11011111100101:	sigmoid_prime = 18'b000001000100110000;
		14'b11011111100110:	sigmoid_prime = 18'b000001000100111000;
		14'b11011111100111:	sigmoid_prime = 18'b000001000101000001;
		14'b11011111101000:	sigmoid_prime = 18'b000001000101001001;
		14'b11011111101001:	sigmoid_prime = 18'b000001000101010001;
		14'b11011111101010:	sigmoid_prime = 18'b000001000101011010;
		14'b11011111101011:	sigmoid_prime = 18'b000001000101100010;
		14'b11011111101100:	sigmoid_prime = 18'b000001000101101010;
		14'b11011111101101:	sigmoid_prime = 18'b000001000101110011;
		14'b11011111101110:	sigmoid_prime = 18'b000001000101111011;
		14'b11011111101111:	sigmoid_prime = 18'b000001000110000100;
		14'b11011111110000:	sigmoid_prime = 18'b000001000110001100;
		14'b11011111110001:	sigmoid_prime = 18'b000001000110010101;
		14'b11011111110010:	sigmoid_prime = 18'b000001000110011101;
		14'b11011111110011:	sigmoid_prime = 18'b000001000110100110;
		14'b11011111110100:	sigmoid_prime = 18'b000001000110101110;
		14'b11011111110101:	sigmoid_prime = 18'b000001000110110111;
		14'b11011111110110:	sigmoid_prime = 18'b000001000110111111;
		14'b11011111110111:	sigmoid_prime = 18'b000001000111001000;
		14'b11011111111000:	sigmoid_prime = 18'b000001000111010000;
		14'b11011111111001:	sigmoid_prime = 18'b000001000111011001;
		14'b11011111111010:	sigmoid_prime = 18'b000001000111100010;
		14'b11011111111011:	sigmoid_prime = 18'b000001000111101010;
		14'b11011111111100:	sigmoid_prime = 18'b000001000111110011;
		14'b11011111111101:	sigmoid_prime = 18'b000001000111111100;
		14'b11011111111110:	sigmoid_prime = 18'b000001001000000100;
		14'b11011111111111:	sigmoid_prime = 18'b000001001000001101;
		14'b11100000000000:	sigmoid_prime = 18'b000001001000010110;
		14'b11100000000001:	sigmoid_prime = 18'b000001001000011110;
		14'b11100000000010:	sigmoid_prime = 18'b000001001000100111;
		14'b11100000000011:	sigmoid_prime = 18'b000001001000110000;
		14'b11100000000100:	sigmoid_prime = 18'b000001001000111001;
		14'b11100000000101:	sigmoid_prime = 18'b000001001001000001;
		14'b11100000000110:	sigmoid_prime = 18'b000001001001001010;
		14'b11100000000111:	sigmoid_prime = 18'b000001001001010011;
		14'b11100000001000:	sigmoid_prime = 18'b000001001001011100;
		14'b11100000001001:	sigmoid_prime = 18'b000001001001100101;
		14'b11100000001010:	sigmoid_prime = 18'b000001001001101110;
		14'b11100000001011:	sigmoid_prime = 18'b000001001001110111;
		14'b11100000001100:	sigmoid_prime = 18'b000001001001111111;
		14'b11100000001101:	sigmoid_prime = 18'b000001001010001000;
		14'b11100000001110:	sigmoid_prime = 18'b000001001010010001;
		14'b11100000001111:	sigmoid_prime = 18'b000001001010011010;
		14'b11100000010000:	sigmoid_prime = 18'b000001001010100011;
		14'b11100000010001:	sigmoid_prime = 18'b000001001010101100;
		14'b11100000010010:	sigmoid_prime = 18'b000001001010110101;
		14'b11100000010011:	sigmoid_prime = 18'b000001001010111110;
		14'b11100000010100:	sigmoid_prime = 18'b000001001011000111;
		14'b11100000010101:	sigmoid_prime = 18'b000001001011010000;
		14'b11100000010110:	sigmoid_prime = 18'b000001001011011001;
		14'b11100000010111:	sigmoid_prime = 18'b000001001011100010;
		14'b11100000011000:	sigmoid_prime = 18'b000001001011101100;
		14'b11100000011001:	sigmoid_prime = 18'b000001001011110101;
		14'b11100000011010:	sigmoid_prime = 18'b000001001011111110;
		14'b11100000011011:	sigmoid_prime = 18'b000001001100000111;
		14'b11100000011100:	sigmoid_prime = 18'b000001001100010000;
		14'b11100000011101:	sigmoid_prime = 18'b000001001100011001;
		14'b11100000011110:	sigmoid_prime = 18'b000001001100100010;
		14'b11100000011111:	sigmoid_prime = 18'b000001001100101100;
		14'b11100000100000:	sigmoid_prime = 18'b000001001100110101;
		14'b11100000100001:	sigmoid_prime = 18'b000001001100111110;
		14'b11100000100010:	sigmoid_prime = 18'b000001001101000111;
		14'b11100000100011:	sigmoid_prime = 18'b000001001101010001;
		14'b11100000100100:	sigmoid_prime = 18'b000001001101011010;
		14'b11100000100101:	sigmoid_prime = 18'b000001001101100011;
		14'b11100000100110:	sigmoid_prime = 18'b000001001101101101;
		14'b11100000100111:	sigmoid_prime = 18'b000001001101110110;
		14'b11100000101000:	sigmoid_prime = 18'b000001001101111111;
		14'b11100000101001:	sigmoid_prime = 18'b000001001110001001;
		14'b11100000101010:	sigmoid_prime = 18'b000001001110010010;
		14'b11100000101011:	sigmoid_prime = 18'b000001001110011011;
		14'b11100000101100:	sigmoid_prime = 18'b000001001110100101;
		14'b11100000101101:	sigmoid_prime = 18'b000001001110101110;
		14'b11100000101110:	sigmoid_prime = 18'b000001001110111000;
		14'b11100000101111:	sigmoid_prime = 18'b000001001111000001;
		14'b11100000110000:	sigmoid_prime = 18'b000001001111001011;
		14'b11100000110001:	sigmoid_prime = 18'b000001001111010100;
		14'b11100000110010:	sigmoid_prime = 18'b000001001111011110;
		14'b11100000110011:	sigmoid_prime = 18'b000001001111100111;
		14'b11100000110100:	sigmoid_prime = 18'b000001001111110001;
		14'b11100000110101:	sigmoid_prime = 18'b000001001111111011;
		14'b11100000110110:	sigmoid_prime = 18'b000001010000000100;
		14'b11100000110111:	sigmoid_prime = 18'b000001010000001110;
		14'b11100000111000:	sigmoid_prime = 18'b000001010000010111;
		14'b11100000111001:	sigmoid_prime = 18'b000001010000100001;
		14'b11100000111010:	sigmoid_prime = 18'b000001010000101011;
		14'b11100000111011:	sigmoid_prime = 18'b000001010000110100;
		14'b11100000111100:	sigmoid_prime = 18'b000001010000111110;
		14'b11100000111101:	sigmoid_prime = 18'b000001010001001000;
		14'b11100000111110:	sigmoid_prime = 18'b000001010001010010;
		14'b11100000111111:	sigmoid_prime = 18'b000001010001011011;
		14'b11100001000000:	sigmoid_prime = 18'b000001010001100101;
		14'b11100001000001:	sigmoid_prime = 18'b000001010001101111;
		14'b11100001000010:	sigmoid_prime = 18'b000001010001111001;
		14'b11100001000011:	sigmoid_prime = 18'b000001010010000011;
		14'b11100001000100:	sigmoid_prime = 18'b000001010010001100;
		14'b11100001000101:	sigmoid_prime = 18'b000001010010010110;
		14'b11100001000110:	sigmoid_prime = 18'b000001010010100000;
		14'b11100001000111:	sigmoid_prime = 18'b000001010010101010;
		14'b11100001001000:	sigmoid_prime = 18'b000001010010110100;
		14'b11100001001001:	sigmoid_prime = 18'b000001010010111110;
		14'b11100001001010:	sigmoid_prime = 18'b000001010011001000;
		14'b11100001001011:	sigmoid_prime = 18'b000001010011010010;
		14'b11100001001100:	sigmoid_prime = 18'b000001010011011100;
		14'b11100001001101:	sigmoid_prime = 18'b000001010011100110;
		14'b11100001001110:	sigmoid_prime = 18'b000001010011110000;
		14'b11100001001111:	sigmoid_prime = 18'b000001010011111010;
		14'b11100001010000:	sigmoid_prime = 18'b000001010100000100;
		14'b11100001010001:	sigmoid_prime = 18'b000001010100001110;
		14'b11100001010010:	sigmoid_prime = 18'b000001010100011000;
		14'b11100001010011:	sigmoid_prime = 18'b000001010100100010;
		14'b11100001010100:	sigmoid_prime = 18'b000001010100101100;
		14'b11100001010101:	sigmoid_prime = 18'b000001010100110111;
		14'b11100001010110:	sigmoid_prime = 18'b000001010101000001;
		14'b11100001010111:	sigmoid_prime = 18'b000001010101001011;
		14'b11100001011000:	sigmoid_prime = 18'b000001010101010101;
		14'b11100001011001:	sigmoid_prime = 18'b000001010101011111;
		14'b11100001011010:	sigmoid_prime = 18'b000001010101101010;
		14'b11100001011011:	sigmoid_prime = 18'b000001010101110100;
		14'b11100001011100:	sigmoid_prime = 18'b000001010101111110;
		14'b11100001011101:	sigmoid_prime = 18'b000001010110001000;
		14'b11100001011110:	sigmoid_prime = 18'b000001010110010011;
		14'b11100001011111:	sigmoid_prime = 18'b000001010110011101;
		14'b11100001100000:	sigmoid_prime = 18'b000001010110100111;
		14'b11100001100001:	sigmoid_prime = 18'b000001010110110010;
		14'b11100001100010:	sigmoid_prime = 18'b000001010110111100;
		14'b11100001100011:	sigmoid_prime = 18'b000001010111000111;
		14'b11100001100100:	sigmoid_prime = 18'b000001010111010001;
		14'b11100001100101:	sigmoid_prime = 18'b000001010111011011;
		14'b11100001100110:	sigmoid_prime = 18'b000001010111100110;
		14'b11100001100111:	sigmoid_prime = 18'b000001010111110000;
		14'b11100001101000:	sigmoid_prime = 18'b000001010111111011;
		14'b11100001101001:	sigmoid_prime = 18'b000001011000000101;
		14'b11100001101010:	sigmoid_prime = 18'b000001011000010000;
		14'b11100001101011:	sigmoid_prime = 18'b000001011000011010;
		14'b11100001101100:	sigmoid_prime = 18'b000001011000100101;
		14'b11100001101101:	sigmoid_prime = 18'b000001011000110000;
		14'b11100001101110:	sigmoid_prime = 18'b000001011000111010;
		14'b11100001101111:	sigmoid_prime = 18'b000001011001000101;
		14'b11100001110000:	sigmoid_prime = 18'b000001011001001111;
		14'b11100001110001:	sigmoid_prime = 18'b000001011001011010;
		14'b11100001110010:	sigmoid_prime = 18'b000001011001100101;
		14'b11100001110011:	sigmoid_prime = 18'b000001011001110000;
		14'b11100001110100:	sigmoid_prime = 18'b000001011001111010;
		14'b11100001110101:	sigmoid_prime = 18'b000001011010000101;
		14'b11100001110110:	sigmoid_prime = 18'b000001011010010000;
		14'b11100001110111:	sigmoid_prime = 18'b000001011010011011;
		14'b11100001111000:	sigmoid_prime = 18'b000001011010100101;
		14'b11100001111001:	sigmoid_prime = 18'b000001011010110000;
		14'b11100001111010:	sigmoid_prime = 18'b000001011010111011;
		14'b11100001111011:	sigmoid_prime = 18'b000001011011000110;
		14'b11100001111100:	sigmoid_prime = 18'b000001011011010001;
		14'b11100001111101:	sigmoid_prime = 18'b000001011011011100;
		14'b11100001111110:	sigmoid_prime = 18'b000001011011100111;
		14'b11100001111111:	sigmoid_prime = 18'b000001011011110010;
		14'b11100010000000:	sigmoid_prime = 18'b000001011011111100;
		14'b11100010000001:	sigmoid_prime = 18'b000001011100000111;
		14'b11100010000010:	sigmoid_prime = 18'b000001011100010010;
		14'b11100010000011:	sigmoid_prime = 18'b000001011100011101;
		14'b11100010000100:	sigmoid_prime = 18'b000001011100101000;
		14'b11100010000101:	sigmoid_prime = 18'b000001011100110100;
		14'b11100010000110:	sigmoid_prime = 18'b000001011100111111;
		14'b11100010000111:	sigmoid_prime = 18'b000001011101001010;
		14'b11100010001000:	sigmoid_prime = 18'b000001011101010101;
		14'b11100010001001:	sigmoid_prime = 18'b000001011101100000;
		14'b11100010001010:	sigmoid_prime = 18'b000001011101101011;
		14'b11100010001011:	sigmoid_prime = 18'b000001011101110110;
		14'b11100010001100:	sigmoid_prime = 18'b000001011110000001;
		14'b11100010001101:	sigmoid_prime = 18'b000001011110001101;
		14'b11100010001110:	sigmoid_prime = 18'b000001011110011000;
		14'b11100010001111:	sigmoid_prime = 18'b000001011110100011;
		14'b11100010010000:	sigmoid_prime = 18'b000001011110101110;
		14'b11100010010001:	sigmoid_prime = 18'b000001011110111010;
		14'b11100010010010:	sigmoid_prime = 18'b000001011111000101;
		14'b11100010010011:	sigmoid_prime = 18'b000001011111010000;
		14'b11100010010100:	sigmoid_prime = 18'b000001011111011100;
		14'b11100010010101:	sigmoid_prime = 18'b000001011111100111;
		14'b11100010010110:	sigmoid_prime = 18'b000001011111110010;
		14'b11100010010111:	sigmoid_prime = 18'b000001011111111110;
		14'b11100010011000:	sigmoid_prime = 18'b000001100000001001;
		14'b11100010011001:	sigmoid_prime = 18'b000001100000010101;
		14'b11100010011010:	sigmoid_prime = 18'b000001100000100000;
		14'b11100010011011:	sigmoid_prime = 18'b000001100000101100;
		14'b11100010011100:	sigmoid_prime = 18'b000001100000110111;
		14'b11100010011101:	sigmoid_prime = 18'b000001100001000011;
		14'b11100010011110:	sigmoid_prime = 18'b000001100001001110;
		14'b11100010011111:	sigmoid_prime = 18'b000001100001011010;
		14'b11100010100000:	sigmoid_prime = 18'b000001100001100110;
		14'b11100010100001:	sigmoid_prime = 18'b000001100001110001;
		14'b11100010100010:	sigmoid_prime = 18'b000001100001111101;
		14'b11100010100011:	sigmoid_prime = 18'b000001100010001000;
		14'b11100010100100:	sigmoid_prime = 18'b000001100010010100;
		14'b11100010100101:	sigmoid_prime = 18'b000001100010100000;
		14'b11100010100110:	sigmoid_prime = 18'b000001100010101011;
		14'b11100010100111:	sigmoid_prime = 18'b000001100010110111;
		14'b11100010101000:	sigmoid_prime = 18'b000001100011000011;
		14'b11100010101001:	sigmoid_prime = 18'b000001100011001111;
		14'b11100010101010:	sigmoid_prime = 18'b000001100011011011;
		14'b11100010101011:	sigmoid_prime = 18'b000001100011100110;
		14'b11100010101100:	sigmoid_prime = 18'b000001100011110010;
		14'b11100010101101:	sigmoid_prime = 18'b000001100011111110;
		14'b11100010101110:	sigmoid_prime = 18'b000001100100001010;
		14'b11100010101111:	sigmoid_prime = 18'b000001100100010110;
		14'b11100010110000:	sigmoid_prime = 18'b000001100100100010;
		14'b11100010110001:	sigmoid_prime = 18'b000001100100101110;
		14'b11100010110010:	sigmoid_prime = 18'b000001100100111010;
		14'b11100010110011:	sigmoid_prime = 18'b000001100101000110;
		14'b11100010110100:	sigmoid_prime = 18'b000001100101010010;
		14'b11100010110101:	sigmoid_prime = 18'b000001100101011110;
		14'b11100010110110:	sigmoid_prime = 18'b000001100101101010;
		14'b11100010110111:	sigmoid_prime = 18'b000001100101110110;
		14'b11100010111000:	sigmoid_prime = 18'b000001100110000010;
		14'b11100010111001:	sigmoid_prime = 18'b000001100110001110;
		14'b11100010111010:	sigmoid_prime = 18'b000001100110011010;
		14'b11100010111011:	sigmoid_prime = 18'b000001100110100110;
		14'b11100010111100:	sigmoid_prime = 18'b000001100110110011;
		14'b11100010111101:	sigmoid_prime = 18'b000001100110111111;
		14'b11100010111110:	sigmoid_prime = 18'b000001100111001011;
		14'b11100010111111:	sigmoid_prime = 18'b000001100111010111;
		14'b11100011000000:	sigmoid_prime = 18'b000001100111100011;
		14'b11100011000001:	sigmoid_prime = 18'b000001100111110000;
		14'b11100011000010:	sigmoid_prime = 18'b000001100111111100;
		14'b11100011000011:	sigmoid_prime = 18'b000001101000001000;
		14'b11100011000100:	sigmoid_prime = 18'b000001101000010101;
		14'b11100011000101:	sigmoid_prime = 18'b000001101000100001;
		14'b11100011000110:	sigmoid_prime = 18'b000001101000101101;
		14'b11100011000111:	sigmoid_prime = 18'b000001101000111010;
		14'b11100011001000:	sigmoid_prime = 18'b000001101001000110;
		14'b11100011001001:	sigmoid_prime = 18'b000001101001010011;
		14'b11100011001010:	sigmoid_prime = 18'b000001101001011111;
		14'b11100011001011:	sigmoid_prime = 18'b000001101001101100;
		14'b11100011001100:	sigmoid_prime = 18'b000001101001111000;
		14'b11100011001101:	sigmoid_prime = 18'b000001101010000101;
		14'b11100011001110:	sigmoid_prime = 18'b000001101010010001;
		14'b11100011001111:	sigmoid_prime = 18'b000001101010011110;
		14'b11100011010000:	sigmoid_prime = 18'b000001101010101011;
		14'b11100011010001:	sigmoid_prime = 18'b000001101010110111;
		14'b11100011010010:	sigmoid_prime = 18'b000001101011000100;
		14'b11100011010011:	sigmoid_prime = 18'b000001101011010001;
		14'b11100011010100:	sigmoid_prime = 18'b000001101011011101;
		14'b11100011010101:	sigmoid_prime = 18'b000001101011101010;
		14'b11100011010110:	sigmoid_prime = 18'b000001101011110111;
		14'b11100011010111:	sigmoid_prime = 18'b000001101100000011;
		14'b11100011011000:	sigmoid_prime = 18'b000001101100010000;
		14'b11100011011001:	sigmoid_prime = 18'b000001101100011101;
		14'b11100011011010:	sigmoid_prime = 18'b000001101100101010;
		14'b11100011011011:	sigmoid_prime = 18'b000001101100110111;
		14'b11100011011100:	sigmoid_prime = 18'b000001101101000100;
		14'b11100011011101:	sigmoid_prime = 18'b000001101101010001;
		14'b11100011011110:	sigmoid_prime = 18'b000001101101011101;
		14'b11100011011111:	sigmoid_prime = 18'b000001101101101010;
		14'b11100011100000:	sigmoid_prime = 18'b000001101101110111;
		14'b11100011100001:	sigmoid_prime = 18'b000001101110000100;
		14'b11100011100010:	sigmoid_prime = 18'b000001101110010001;
		14'b11100011100011:	sigmoid_prime = 18'b000001101110011110;
		14'b11100011100100:	sigmoid_prime = 18'b000001101110101011;
		14'b11100011100101:	sigmoid_prime = 18'b000001101110111001;
		14'b11100011100110:	sigmoid_prime = 18'b000001101111000110;
		14'b11100011100111:	sigmoid_prime = 18'b000001101111010011;
		14'b11100011101000:	sigmoid_prime = 18'b000001101111100000;
		14'b11100011101001:	sigmoid_prime = 18'b000001101111101101;
		14'b11100011101010:	sigmoid_prime = 18'b000001101111111010;
		14'b11100011101011:	sigmoid_prime = 18'b000001110000000111;
		14'b11100011101100:	sigmoid_prime = 18'b000001110000010101;
		14'b11100011101101:	sigmoid_prime = 18'b000001110000100010;
		14'b11100011101110:	sigmoid_prime = 18'b000001110000101111;
		14'b11100011101111:	sigmoid_prime = 18'b000001110000111101;
		14'b11100011110000:	sigmoid_prime = 18'b000001110001001010;
		14'b11100011110001:	sigmoid_prime = 18'b000001110001010111;
		14'b11100011110010:	sigmoid_prime = 18'b000001110001100101;
		14'b11100011110011:	sigmoid_prime = 18'b000001110001110010;
		14'b11100011110100:	sigmoid_prime = 18'b000001110001111111;
		14'b11100011110101:	sigmoid_prime = 18'b000001110010001101;
		14'b11100011110110:	sigmoid_prime = 18'b000001110010011010;
		14'b11100011110111:	sigmoid_prime = 18'b000001110010101000;
		14'b11100011111000:	sigmoid_prime = 18'b000001110010110101;
		14'b11100011111001:	sigmoid_prime = 18'b000001110011000011;
		14'b11100011111010:	sigmoid_prime = 18'b000001110011010000;
		14'b11100011111011:	sigmoid_prime = 18'b000001110011011110;
		14'b11100011111100:	sigmoid_prime = 18'b000001110011101100;
		14'b11100011111101:	sigmoid_prime = 18'b000001110011111001;
		14'b11100011111110:	sigmoid_prime = 18'b000001110100000111;
		14'b11100011111111:	sigmoid_prime = 18'b000001110100010101;
		14'b11100100000000:	sigmoid_prime = 18'b000001110100100010;
		14'b11100100000001:	sigmoid_prime = 18'b000001110100110000;
		14'b11100100000010:	sigmoid_prime = 18'b000001110100111110;
		14'b11100100000011:	sigmoid_prime = 18'b000001110101001100;
		14'b11100100000100:	sigmoid_prime = 18'b000001110101011001;
		14'b11100100000101:	sigmoid_prime = 18'b000001110101100111;
		14'b11100100000110:	sigmoid_prime = 18'b000001110101110101;
		14'b11100100000111:	sigmoid_prime = 18'b000001110110000011;
		14'b11100100001000:	sigmoid_prime = 18'b000001110110010001;
		14'b11100100001001:	sigmoid_prime = 18'b000001110110011111;
		14'b11100100001010:	sigmoid_prime = 18'b000001110110101101;
		14'b11100100001011:	sigmoid_prime = 18'b000001110110111011;
		14'b11100100001100:	sigmoid_prime = 18'b000001110111001001;
		14'b11100100001101:	sigmoid_prime = 18'b000001110111010111;
		14'b11100100001110:	sigmoid_prime = 18'b000001110111100101;
		14'b11100100001111:	sigmoid_prime = 18'b000001110111110011;
		14'b11100100010000:	sigmoid_prime = 18'b000001111000000001;
		14'b11100100010001:	sigmoid_prime = 18'b000001111000001111;
		14'b11100100010010:	sigmoid_prime = 18'b000001111000011101;
		14'b11100100010011:	sigmoid_prime = 18'b000001111000101011;
		14'b11100100010100:	sigmoid_prime = 18'b000001111000111001;
		14'b11100100010101:	sigmoid_prime = 18'b000001111001001000;
		14'b11100100010110:	sigmoid_prime = 18'b000001111001010110;
		14'b11100100010111:	sigmoid_prime = 18'b000001111001100100;
		14'b11100100011000:	sigmoid_prime = 18'b000001111001110010;
		14'b11100100011001:	sigmoid_prime = 18'b000001111010000001;
		14'b11100100011010:	sigmoid_prime = 18'b000001111010001111;
		14'b11100100011011:	sigmoid_prime = 18'b000001111010011101;
		14'b11100100011100:	sigmoid_prime = 18'b000001111010101100;
		14'b11100100011101:	sigmoid_prime = 18'b000001111010111010;
		14'b11100100011110:	sigmoid_prime = 18'b000001111011001000;
		14'b11100100011111:	sigmoid_prime = 18'b000001111011010111;
		14'b11100100100000:	sigmoid_prime = 18'b000001111011100101;
		14'b11100100100001:	sigmoid_prime = 18'b000001111011110100;
		14'b11100100100010:	sigmoid_prime = 18'b000001111100000010;
		14'b11100100100011:	sigmoid_prime = 18'b000001111100010001;
		14'b11100100100100:	sigmoid_prime = 18'b000001111100100000;
		14'b11100100100101:	sigmoid_prime = 18'b000001111100101110;
		14'b11100100100110:	sigmoid_prime = 18'b000001111100111101;
		14'b11100100100111:	sigmoid_prime = 18'b000001111101001011;
		14'b11100100101000:	sigmoid_prime = 18'b000001111101011010;
		14'b11100100101001:	sigmoid_prime = 18'b000001111101101001;
		14'b11100100101010:	sigmoid_prime = 18'b000001111101111000;
		14'b11100100101011:	sigmoid_prime = 18'b000001111110000110;
		14'b11100100101100:	sigmoid_prime = 18'b000001111110010101;
		14'b11100100101101:	sigmoid_prime = 18'b000001111110100100;
		14'b11100100101110:	sigmoid_prime = 18'b000001111110110011;
		14'b11100100101111:	sigmoid_prime = 18'b000001111111000010;
		14'b11100100110000:	sigmoid_prime = 18'b000001111111010000;
		14'b11100100110001:	sigmoid_prime = 18'b000001111111011111;
		14'b11100100110010:	sigmoid_prime = 18'b000001111111101110;
		14'b11100100110011:	sigmoid_prime = 18'b000001111111111101;
		14'b11100100110100:	sigmoid_prime = 18'b000010000000001100;
		14'b11100100110101:	sigmoid_prime = 18'b000010000000011011;
		14'b11100100110110:	sigmoid_prime = 18'b000010000000101010;
		14'b11100100110111:	sigmoid_prime = 18'b000010000000111001;
		14'b11100100111000:	sigmoid_prime = 18'b000010000001001000;
		14'b11100100111001:	sigmoid_prime = 18'b000010000001010111;
		14'b11100100111010:	sigmoid_prime = 18'b000010000001100111;
		14'b11100100111011:	sigmoid_prime = 18'b000010000001110110;
		14'b11100100111100:	sigmoid_prime = 18'b000010000010000101;
		14'b11100100111101:	sigmoid_prime = 18'b000010000010010100;
		14'b11100100111110:	sigmoid_prime = 18'b000010000010100011;
		14'b11100100111111:	sigmoid_prime = 18'b000010000010110011;
		14'b11100101000000:	sigmoid_prime = 18'b000010000011000010;
		14'b11100101000001:	sigmoid_prime = 18'b000010000011010001;
		14'b11100101000010:	sigmoid_prime = 18'b000010000011100000;
		14'b11100101000011:	sigmoid_prime = 18'b000010000011110000;
		14'b11100101000100:	sigmoid_prime = 18'b000010000011111111;
		14'b11100101000101:	sigmoid_prime = 18'b000010000100001111;
		14'b11100101000110:	sigmoid_prime = 18'b000010000100011110;
		14'b11100101000111:	sigmoid_prime = 18'b000010000100101110;
		14'b11100101001000:	sigmoid_prime = 18'b000010000100111101;
		14'b11100101001001:	sigmoid_prime = 18'b000010000101001101;
		14'b11100101001010:	sigmoid_prime = 18'b000010000101011100;
		14'b11100101001011:	sigmoid_prime = 18'b000010000101101100;
		14'b11100101001100:	sigmoid_prime = 18'b000010000101111011;
		14'b11100101001101:	sigmoid_prime = 18'b000010000110001011;
		14'b11100101001110:	sigmoid_prime = 18'b000010000110011011;
		14'b11100101001111:	sigmoid_prime = 18'b000010000110101010;
		14'b11100101010000:	sigmoid_prime = 18'b000010000110111010;
		14'b11100101010001:	sigmoid_prime = 18'b000010000111001010;
		14'b11100101010010:	sigmoid_prime = 18'b000010000111011001;
		14'b11100101010011:	sigmoid_prime = 18'b000010000111101001;
		14'b11100101010100:	sigmoid_prime = 18'b000010000111111001;
		14'b11100101010101:	sigmoid_prime = 18'b000010001000001001;
		14'b11100101010110:	sigmoid_prime = 18'b000010001000011001;
		14'b11100101010111:	sigmoid_prime = 18'b000010001000101001;
		14'b11100101011000:	sigmoid_prime = 18'b000010001000111000;
		14'b11100101011001:	sigmoid_prime = 18'b000010001001001000;
		14'b11100101011010:	sigmoid_prime = 18'b000010001001011000;
		14'b11100101011011:	sigmoid_prime = 18'b000010001001101000;
		14'b11100101011100:	sigmoid_prime = 18'b000010001001111000;
		14'b11100101011101:	sigmoid_prime = 18'b000010001010001000;
		14'b11100101011110:	sigmoid_prime = 18'b000010001010011000;
		14'b11100101011111:	sigmoid_prime = 18'b000010001010101001;
		14'b11100101100000:	sigmoid_prime = 18'b000010001010111001;
		14'b11100101100001:	sigmoid_prime = 18'b000010001011001001;
		14'b11100101100010:	sigmoid_prime = 18'b000010001011011001;
		14'b11100101100011:	sigmoid_prime = 18'b000010001011101001;
		14'b11100101100100:	sigmoid_prime = 18'b000010001011111010;
		14'b11100101100101:	sigmoid_prime = 18'b000010001100001010;
		14'b11100101100110:	sigmoid_prime = 18'b000010001100011010;
		14'b11100101100111:	sigmoid_prime = 18'b000010001100101010;
		14'b11100101101000:	sigmoid_prime = 18'b000010001100111011;
		14'b11100101101001:	sigmoid_prime = 18'b000010001101001011;
		14'b11100101101010:	sigmoid_prime = 18'b000010001101011011;
		14'b11100101101011:	sigmoid_prime = 18'b000010001101101100;
		14'b11100101101100:	sigmoid_prime = 18'b000010001101111100;
		14'b11100101101101:	sigmoid_prime = 18'b000010001110001101;
		14'b11100101101110:	sigmoid_prime = 18'b000010001110011101;
		14'b11100101101111:	sigmoid_prime = 18'b000010001110101110;
		14'b11100101110000:	sigmoid_prime = 18'b000010001110111110;
		14'b11100101110001:	sigmoid_prime = 18'b000010001111001111;
		14'b11100101110010:	sigmoid_prime = 18'b000010001111100000;
		14'b11100101110011:	sigmoid_prime = 18'b000010001111110000;
		14'b11100101110100:	sigmoid_prime = 18'b000010010000000001;
		14'b11100101110101:	sigmoid_prime = 18'b000010010000010010;
		14'b11100101110110:	sigmoid_prime = 18'b000010010000100010;
		14'b11100101110111:	sigmoid_prime = 18'b000010010000110011;
		14'b11100101111000:	sigmoid_prime = 18'b000010010001000100;
		14'b11100101111001:	sigmoid_prime = 18'b000010010001010101;
		14'b11100101111010:	sigmoid_prime = 18'b000010010001100110;
		14'b11100101111011:	sigmoid_prime = 18'b000010010001110111;
		14'b11100101111100:	sigmoid_prime = 18'b000010010010000111;
		14'b11100101111101:	sigmoid_prime = 18'b000010010010011000;
		14'b11100101111110:	sigmoid_prime = 18'b000010010010101001;
		14'b11100101111111:	sigmoid_prime = 18'b000010010010111010;
		14'b11100110000000:	sigmoid_prime = 18'b000010010011001011;
		14'b11100110000001:	sigmoid_prime = 18'b000010010011011100;
		14'b11100110000010:	sigmoid_prime = 18'b000010010011101101;
		14'b11100110000011:	sigmoid_prime = 18'b000010010011111110;
		14'b11100110000100:	sigmoid_prime = 18'b000010010100010000;
		14'b11100110000101:	sigmoid_prime = 18'b000010010100100001;
		14'b11100110000110:	sigmoid_prime = 18'b000010010100110010;
		14'b11100110000111:	sigmoid_prime = 18'b000010010101000011;
		14'b11100110001000:	sigmoid_prime = 18'b000010010101010100;
		14'b11100110001001:	sigmoid_prime = 18'b000010010101100110;
		14'b11100110001010:	sigmoid_prime = 18'b000010010101110111;
		14'b11100110001011:	sigmoid_prime = 18'b000010010110001000;
		14'b11100110001100:	sigmoid_prime = 18'b000010010110011010;
		14'b11100110001101:	sigmoid_prime = 18'b000010010110101011;
		14'b11100110001110:	sigmoid_prime = 18'b000010010110111100;
		14'b11100110001111:	sigmoid_prime = 18'b000010010111001110;
		14'b11100110010000:	sigmoid_prime = 18'b000010010111011111;
		14'b11100110010001:	sigmoid_prime = 18'b000010010111110001;
		14'b11100110010010:	sigmoid_prime = 18'b000010011000000010;
		14'b11100110010011:	sigmoid_prime = 18'b000010011000010100;
		14'b11100110010100:	sigmoid_prime = 18'b000010011000100101;
		14'b11100110010101:	sigmoid_prime = 18'b000010011000110111;
		14'b11100110010110:	sigmoid_prime = 18'b000010011001001001;
		14'b11100110010111:	sigmoid_prime = 18'b000010011001011010;
		14'b11100110011000:	sigmoid_prime = 18'b000010011001101100;
		14'b11100110011001:	sigmoid_prime = 18'b000010011001111110;
		14'b11100110011010:	sigmoid_prime = 18'b000010011010010000;
		14'b11100110011011:	sigmoid_prime = 18'b000010011010100001;
		14'b11100110011100:	sigmoid_prime = 18'b000010011010110011;
		14'b11100110011101:	sigmoid_prime = 18'b000010011011000101;
		14'b11100110011110:	sigmoid_prime = 18'b000010011011010111;
		14'b11100110011111:	sigmoid_prime = 18'b000010011011101001;
		14'b11100110100000:	sigmoid_prime = 18'b000010011011111011;
		14'b11100110100001:	sigmoid_prime = 18'b000010011100001101;
		14'b11100110100010:	sigmoid_prime = 18'b000010011100011111;
		14'b11100110100011:	sigmoid_prime = 18'b000010011100110001;
		14'b11100110100100:	sigmoid_prime = 18'b000010011101000011;
		14'b11100110100101:	sigmoid_prime = 18'b000010011101010101;
		14'b11100110100110:	sigmoid_prime = 18'b000010011101100111;
		14'b11100110100111:	sigmoid_prime = 18'b000010011101111001;
		14'b11100110101000:	sigmoid_prime = 18'b000010011110001011;
		14'b11100110101001:	sigmoid_prime = 18'b000010011110011101;
		14'b11100110101010:	sigmoid_prime = 18'b000010011110110000;
		14'b11100110101011:	sigmoid_prime = 18'b000010011111000010;
		14'b11100110101100:	sigmoid_prime = 18'b000010011111010100;
		14'b11100110101101:	sigmoid_prime = 18'b000010011111100110;
		14'b11100110101110:	sigmoid_prime = 18'b000010011111111001;
		14'b11100110101111:	sigmoid_prime = 18'b000010100000001011;
		14'b11100110110000:	sigmoid_prime = 18'b000010100000011110;
		14'b11100110110001:	sigmoid_prime = 18'b000010100000110000;
		14'b11100110110010:	sigmoid_prime = 18'b000010100001000011;
		14'b11100110110011:	sigmoid_prime = 18'b000010100001010101;
		14'b11100110110100:	sigmoid_prime = 18'b000010100001101000;
		14'b11100110110101:	sigmoid_prime = 18'b000010100001111010;
		14'b11100110110110:	sigmoid_prime = 18'b000010100010001101;
		14'b11100110110111:	sigmoid_prime = 18'b000010100010011111;
		14'b11100110111000:	sigmoid_prime = 18'b000010100010110010;
		14'b11100110111001:	sigmoid_prime = 18'b000010100011000101;
		14'b11100110111010:	sigmoid_prime = 18'b000010100011010111;
		14'b11100110111011:	sigmoid_prime = 18'b000010100011101010;
		14'b11100110111100:	sigmoid_prime = 18'b000010100011111101;
		14'b11100110111101:	sigmoid_prime = 18'b000010100100010000;
		14'b11100110111110:	sigmoid_prime = 18'b000010100100100010;
		14'b11100110111111:	sigmoid_prime = 18'b000010100100110101;
		14'b11100111000000:	sigmoid_prime = 18'b000010100101001000;
		14'b11100111000001:	sigmoid_prime = 18'b000010100101011011;
		14'b11100111000010:	sigmoid_prime = 18'b000010100101101110;
		14'b11100111000011:	sigmoid_prime = 18'b000010100110000001;
		14'b11100111000100:	sigmoid_prime = 18'b000010100110010100;
		14'b11100111000101:	sigmoid_prime = 18'b000010100110100111;
		14'b11100111000110:	sigmoid_prime = 18'b000010100110111010;
		14'b11100111000111:	sigmoid_prime = 18'b000010100111001101;
		14'b11100111001000:	sigmoid_prime = 18'b000010100111100000;
		14'b11100111001001:	sigmoid_prime = 18'b000010100111110100;
		14'b11100111001010:	sigmoid_prime = 18'b000010101000000111;
		14'b11100111001011:	sigmoid_prime = 18'b000010101000011010;
		14'b11100111001100:	sigmoid_prime = 18'b000010101000101101;
		14'b11100111001101:	sigmoid_prime = 18'b000010101001000001;
		14'b11100111001110:	sigmoid_prime = 18'b000010101001010100;
		14'b11100111001111:	sigmoid_prime = 18'b000010101001100111;
		14'b11100111010000:	sigmoid_prime = 18'b000010101001111011;
		14'b11100111010001:	sigmoid_prime = 18'b000010101010001110;
		14'b11100111010010:	sigmoid_prime = 18'b000010101010100001;
		14'b11100111010011:	sigmoid_prime = 18'b000010101010110101;
		14'b11100111010100:	sigmoid_prime = 18'b000010101011001000;
		14'b11100111010101:	sigmoid_prime = 18'b000010101011011100;
		14'b11100111010110:	sigmoid_prime = 18'b000010101011110000;
		14'b11100111010111:	sigmoid_prime = 18'b000010101100000011;
		14'b11100111011000:	sigmoid_prime = 18'b000010101100010111;
		14'b11100111011001:	sigmoid_prime = 18'b000010101100101010;
		14'b11100111011010:	sigmoid_prime = 18'b000010101100111110;
		14'b11100111011011:	sigmoid_prime = 18'b000010101101010010;
		14'b11100111011100:	sigmoid_prime = 18'b000010101101100110;
		14'b11100111011101:	sigmoid_prime = 18'b000010101101111001;
		14'b11100111011110:	sigmoid_prime = 18'b000010101110001101;
		14'b11100111011111:	sigmoid_prime = 18'b000010101110100001;
		14'b11100111100000:	sigmoid_prime = 18'b000010101110110101;
		14'b11100111100001:	sigmoid_prime = 18'b000010101111001001;
		14'b11100111100010:	sigmoid_prime = 18'b000010101111011101;
		14'b11100111100011:	sigmoid_prime = 18'b000010101111110001;
		14'b11100111100100:	sigmoid_prime = 18'b000010110000000101;
		14'b11100111100101:	sigmoid_prime = 18'b000010110000011001;
		14'b11100111100110:	sigmoid_prime = 18'b000010110000101101;
		14'b11100111100111:	sigmoid_prime = 18'b000010110001000001;
		14'b11100111101000:	sigmoid_prime = 18'b000010110001010101;
		14'b11100111101001:	sigmoid_prime = 18'b000010110001101001;
		14'b11100111101010:	sigmoid_prime = 18'b000010110001111110;
		14'b11100111101011:	sigmoid_prime = 18'b000010110010010010;
		14'b11100111101100:	sigmoid_prime = 18'b000010110010100110;
		14'b11100111101101:	sigmoid_prime = 18'b000010110010111010;
		14'b11100111101110:	sigmoid_prime = 18'b000010110011001111;
		14'b11100111101111:	sigmoid_prime = 18'b000010110011100011;
		14'b11100111110000:	sigmoid_prime = 18'b000010110011110111;
		14'b11100111110001:	sigmoid_prime = 18'b000010110100001100;
		14'b11100111110010:	sigmoid_prime = 18'b000010110100100000;
		14'b11100111110011:	sigmoid_prime = 18'b000010110100110101;
		14'b11100111110100:	sigmoid_prime = 18'b000010110101001001;
		14'b11100111110101:	sigmoid_prime = 18'b000010110101011110;
		14'b11100111110110:	sigmoid_prime = 18'b000010110101110011;
		14'b11100111110111:	sigmoid_prime = 18'b000010110110000111;
		14'b11100111111000:	sigmoid_prime = 18'b000010110110011100;
		14'b11100111111001:	sigmoid_prime = 18'b000010110110110001;
		14'b11100111111010:	sigmoid_prime = 18'b000010110111000101;
		14'b11100111111011:	sigmoid_prime = 18'b000010110111011010;
		14'b11100111111100:	sigmoid_prime = 18'b000010110111101111;
		14'b11100111111101:	sigmoid_prime = 18'b000010111000000100;
		14'b11100111111110:	sigmoid_prime = 18'b000010111000011000;
		14'b11100111111111:	sigmoid_prime = 18'b000010111000101101;
		14'b11101000000000:	sigmoid_prime = 18'b000010111001000010;
		14'b11101000000001:	sigmoid_prime = 18'b000010111001010111;
		14'b11101000000010:	sigmoid_prime = 18'b000010111001101100;
		14'b11101000000011:	sigmoid_prime = 18'b000010111010000001;
		14'b11101000000100:	sigmoid_prime = 18'b000010111010010110;
		14'b11101000000101:	sigmoid_prime = 18'b000010111010101011;
		14'b11101000000110:	sigmoid_prime = 18'b000010111011000001;
		14'b11101000000111:	sigmoid_prime = 18'b000010111011010110;
		14'b11101000001000:	sigmoid_prime = 18'b000010111011101011;
		14'b11101000001001:	sigmoid_prime = 18'b000010111100000000;
		14'b11101000001010:	sigmoid_prime = 18'b000010111100010101;
		14'b11101000001011:	sigmoid_prime = 18'b000010111100101011;
		14'b11101000001100:	sigmoid_prime = 18'b000010111101000000;
		14'b11101000001101:	sigmoid_prime = 18'b000010111101010101;
		14'b11101000001110:	sigmoid_prime = 18'b000010111101101011;
		14'b11101000001111:	sigmoid_prime = 18'b000010111110000000;
		14'b11101000010000:	sigmoid_prime = 18'b000010111110010110;
		14'b11101000010001:	sigmoid_prime = 18'b000010111110101011;
		14'b11101000010010:	sigmoid_prime = 18'b000010111111000001;
		14'b11101000010011:	sigmoid_prime = 18'b000010111111010110;
		14'b11101000010100:	sigmoid_prime = 18'b000010111111101100;
		14'b11101000010101:	sigmoid_prime = 18'b000011000000000001;
		14'b11101000010110:	sigmoid_prime = 18'b000011000000010111;
		14'b11101000010111:	sigmoid_prime = 18'b000011000000101101;
		14'b11101000011000:	sigmoid_prime = 18'b000011000001000010;
		14'b11101000011001:	sigmoid_prime = 18'b000011000001011000;
		14'b11101000011010:	sigmoid_prime = 18'b000011000001101110;
		14'b11101000011011:	sigmoid_prime = 18'b000011000010000100;
		14'b11101000011100:	sigmoid_prime = 18'b000011000010011010;
		14'b11101000011101:	sigmoid_prime = 18'b000011000010101111;
		14'b11101000011110:	sigmoid_prime = 18'b000011000011000101;
		14'b11101000011111:	sigmoid_prime = 18'b000011000011011011;
		14'b11101000100000:	sigmoid_prime = 18'b000011000011110001;
		14'b11101000100001:	sigmoid_prime = 18'b000011000100000111;
		14'b11101000100010:	sigmoid_prime = 18'b000011000100011101;
		14'b11101000100011:	sigmoid_prime = 18'b000011000100110011;
		14'b11101000100100:	sigmoid_prime = 18'b000011000101001010;
		14'b11101000100101:	sigmoid_prime = 18'b000011000101100000;
		14'b11101000100110:	sigmoid_prime = 18'b000011000101110110;
		14'b11101000100111:	sigmoid_prime = 18'b000011000110001100;
		14'b11101000101000:	sigmoid_prime = 18'b000011000110100010;
		14'b11101000101001:	sigmoid_prime = 18'b000011000110111001;
		14'b11101000101010:	sigmoid_prime = 18'b000011000111001111;
		14'b11101000101011:	sigmoid_prime = 18'b000011000111100101;
		14'b11101000101100:	sigmoid_prime = 18'b000011000111111100;
		14'b11101000101101:	sigmoid_prime = 18'b000011001000010010;
		14'b11101000101110:	sigmoid_prime = 18'b000011001000101001;
		14'b11101000101111:	sigmoid_prime = 18'b000011001000111111;
		14'b11101000110000:	sigmoid_prime = 18'b000011001001010110;
		14'b11101000110001:	sigmoid_prime = 18'b000011001001101100;
		14'b11101000110010:	sigmoid_prime = 18'b000011001010000011;
		14'b11101000110011:	sigmoid_prime = 18'b000011001010011010;
		14'b11101000110100:	sigmoid_prime = 18'b000011001010110000;
		14'b11101000110101:	sigmoid_prime = 18'b000011001011000111;
		14'b11101000110110:	sigmoid_prime = 18'b000011001011011110;
		14'b11101000110111:	sigmoid_prime = 18'b000011001011110101;
		14'b11101000111000:	sigmoid_prime = 18'b000011001100001011;
		14'b11101000111001:	sigmoid_prime = 18'b000011001100100010;
		14'b11101000111010:	sigmoid_prime = 18'b000011001100111001;
		14'b11101000111011:	sigmoid_prime = 18'b000011001101010000;
		14'b11101000111100:	sigmoid_prime = 18'b000011001101100111;
		14'b11101000111101:	sigmoid_prime = 18'b000011001101111110;
		14'b11101000111110:	sigmoid_prime = 18'b000011001110010101;
		14'b11101000111111:	sigmoid_prime = 18'b000011001110101100;
		14'b11101001000000:	sigmoid_prime = 18'b000011001111000011;
		14'b11101001000001:	sigmoid_prime = 18'b000011001111011010;
		14'b11101001000010:	sigmoid_prime = 18'b000011001111110010;
		14'b11101001000011:	sigmoid_prime = 18'b000011010000001001;
		14'b11101001000100:	sigmoid_prime = 18'b000011010000100000;
		14'b11101001000101:	sigmoid_prime = 18'b000011010000110111;
		14'b11101001000110:	sigmoid_prime = 18'b000011010001001111;
		14'b11101001000111:	sigmoid_prime = 18'b000011010001100110;
		14'b11101001001000:	sigmoid_prime = 18'b000011010001111101;
		14'b11101001001001:	sigmoid_prime = 18'b000011010010010101;
		14'b11101001001010:	sigmoid_prime = 18'b000011010010101100;
		14'b11101001001011:	sigmoid_prime = 18'b000011010011000100;
		14'b11101001001100:	sigmoid_prime = 18'b000011010011011011;
		14'b11101001001101:	sigmoid_prime = 18'b000011010011110011;
		14'b11101001001110:	sigmoid_prime = 18'b000011010100001010;
		14'b11101001001111:	sigmoid_prime = 18'b000011010100100010;
		14'b11101001010000:	sigmoid_prime = 18'b000011010100111010;
		14'b11101001010001:	sigmoid_prime = 18'b000011010101010001;
		14'b11101001010010:	sigmoid_prime = 18'b000011010101101001;
		14'b11101001010011:	sigmoid_prime = 18'b000011010110000001;
		14'b11101001010100:	sigmoid_prime = 18'b000011010110011001;
		14'b11101001010101:	sigmoid_prime = 18'b000011010110110001;
		14'b11101001010110:	sigmoid_prime = 18'b000011010111001000;
		14'b11101001010111:	sigmoid_prime = 18'b000011010111100000;
		14'b11101001011000:	sigmoid_prime = 18'b000011010111111000;
		14'b11101001011001:	sigmoid_prime = 18'b000011011000010000;
		14'b11101001011010:	sigmoid_prime = 18'b000011011000101000;
		14'b11101001011011:	sigmoid_prime = 18'b000011011001000000;
		14'b11101001011100:	sigmoid_prime = 18'b000011011001011000;
		14'b11101001011101:	sigmoid_prime = 18'b000011011001110001;
		14'b11101001011110:	sigmoid_prime = 18'b000011011010001001;
		14'b11101001011111:	sigmoid_prime = 18'b000011011010100001;
		14'b11101001100000:	sigmoid_prime = 18'b000011011010111001;
		14'b11101001100001:	sigmoid_prime = 18'b000011011011010010;
		14'b11101001100010:	sigmoid_prime = 18'b000011011011101010;
		14'b11101001100011:	sigmoid_prime = 18'b000011011100000010;
		14'b11101001100100:	sigmoid_prime = 18'b000011011100011011;
		14'b11101001100101:	sigmoid_prime = 18'b000011011100110011;
		14'b11101001100110:	sigmoid_prime = 18'b000011011101001011;
		14'b11101001100111:	sigmoid_prime = 18'b000011011101100100;
		14'b11101001101000:	sigmoid_prime = 18'b000011011101111101;
		14'b11101001101001:	sigmoid_prime = 18'b000011011110010101;
		14'b11101001101010:	sigmoid_prime = 18'b000011011110101110;
		14'b11101001101011:	sigmoid_prime = 18'b000011011111000110;
		14'b11101001101100:	sigmoid_prime = 18'b000011011111011111;
		14'b11101001101101:	sigmoid_prime = 18'b000011011111111000;
		14'b11101001101110:	sigmoid_prime = 18'b000011100000010000;
		14'b11101001101111:	sigmoid_prime = 18'b000011100000101001;
		14'b11101001110000:	sigmoid_prime = 18'b000011100001000010;
		14'b11101001110001:	sigmoid_prime = 18'b000011100001011011;
		14'b11101001110010:	sigmoid_prime = 18'b000011100001110100;
		14'b11101001110011:	sigmoid_prime = 18'b000011100010001101;
		14'b11101001110100:	sigmoid_prime = 18'b000011100010100110;
		14'b11101001110101:	sigmoid_prime = 18'b000011100010111111;
		14'b11101001110110:	sigmoid_prime = 18'b000011100011011000;
		14'b11101001110111:	sigmoid_prime = 18'b000011100011110001;
		14'b11101001111000:	sigmoid_prime = 18'b000011100100001010;
		14'b11101001111001:	sigmoid_prime = 18'b000011100100100011;
		14'b11101001111010:	sigmoid_prime = 18'b000011100100111100;
		14'b11101001111011:	sigmoid_prime = 18'b000011100101010110;
		14'b11101001111100:	sigmoid_prime = 18'b000011100101101111;
		14'b11101001111101:	sigmoid_prime = 18'b000011100110001000;
		14'b11101001111110:	sigmoid_prime = 18'b000011100110100010;
		14'b11101001111111:	sigmoid_prime = 18'b000011100110111011;
		14'b11101010000000:	sigmoid_prime = 18'b000011100111010100;
		14'b11101010000001:	sigmoid_prime = 18'b000011100111101110;
		14'b11101010000010:	sigmoid_prime = 18'b000011101000000111;
		14'b11101010000011:	sigmoid_prime = 18'b000011101000100001;
		14'b11101010000100:	sigmoid_prime = 18'b000011101000111010;
		14'b11101010000101:	sigmoid_prime = 18'b000011101001010100;
		14'b11101010000110:	sigmoid_prime = 18'b000011101001101110;
		14'b11101010000111:	sigmoid_prime = 18'b000011101010000111;
		14'b11101010001000:	sigmoid_prime = 18'b000011101010100001;
		14'b11101010001001:	sigmoid_prime = 18'b000011101010111011;
		14'b11101010001010:	sigmoid_prime = 18'b000011101011010101;
		14'b11101010001011:	sigmoid_prime = 18'b000011101011101111;
		14'b11101010001100:	sigmoid_prime = 18'b000011101100001000;
		14'b11101010001101:	sigmoid_prime = 18'b000011101100100010;
		14'b11101010001110:	sigmoid_prime = 18'b000011101100111100;
		14'b11101010001111:	sigmoid_prime = 18'b000011101101010110;
		14'b11101010010000:	sigmoid_prime = 18'b000011101101110000;
		14'b11101010010001:	sigmoid_prime = 18'b000011101110001010;
		14'b11101010010010:	sigmoid_prime = 18'b000011101110100100;
		14'b11101010010011:	sigmoid_prime = 18'b000011101110111111;
		14'b11101010010100:	sigmoid_prime = 18'b000011101111011001;
		14'b11101010010101:	sigmoid_prime = 18'b000011101111110011;
		14'b11101010010110:	sigmoid_prime = 18'b000011110000001101;
		14'b11101010010111:	sigmoid_prime = 18'b000011110000100111;
		14'b11101010011000:	sigmoid_prime = 18'b000011110001000010;
		14'b11101010011001:	sigmoid_prime = 18'b000011110001011100;
		14'b11101010011010:	sigmoid_prime = 18'b000011110001110111;
		14'b11101010011011:	sigmoid_prime = 18'b000011110010010001;
		14'b11101010011100:	sigmoid_prime = 18'b000011110010101100;
		14'b11101010011101:	sigmoid_prime = 18'b000011110011000110;
		14'b11101010011110:	sigmoid_prime = 18'b000011110011100001;
		14'b11101010011111:	sigmoid_prime = 18'b000011110011111011;
		14'b11101010100000:	sigmoid_prime = 18'b000011110100010110;
		14'b11101010100001:	sigmoid_prime = 18'b000011110100110000;
		14'b11101010100010:	sigmoid_prime = 18'b000011110101001011;
		14'b11101010100011:	sigmoid_prime = 18'b000011110101100110;
		14'b11101010100100:	sigmoid_prime = 18'b000011110110000001;
		14'b11101010100101:	sigmoid_prime = 18'b000011110110011100;
		14'b11101010100110:	sigmoid_prime = 18'b000011110110110110;
		14'b11101010100111:	sigmoid_prime = 18'b000011110111010001;
		14'b11101010101000:	sigmoid_prime = 18'b000011110111101100;
		14'b11101010101001:	sigmoid_prime = 18'b000011111000000111;
		14'b11101010101010:	sigmoid_prime = 18'b000011111000100010;
		14'b11101010101011:	sigmoid_prime = 18'b000011111000111101;
		14'b11101010101100:	sigmoid_prime = 18'b000011111001011000;
		14'b11101010101101:	sigmoid_prime = 18'b000011111001110100;
		14'b11101010101110:	sigmoid_prime = 18'b000011111010001111;
		14'b11101010101111:	sigmoid_prime = 18'b000011111010101010;
		14'b11101010110000:	sigmoid_prime = 18'b000011111011000101;
		14'b11101010110001:	sigmoid_prime = 18'b000011111011100000;
		14'b11101010110010:	sigmoid_prime = 18'b000011111011111100;
		14'b11101010110011:	sigmoid_prime = 18'b000011111100010111;
		14'b11101010110100:	sigmoid_prime = 18'b000011111100110011;
		14'b11101010110101:	sigmoid_prime = 18'b000011111101001110;
		14'b11101010110110:	sigmoid_prime = 18'b000011111101101001;
		14'b11101010110111:	sigmoid_prime = 18'b000011111110000101;
		14'b11101010111000:	sigmoid_prime = 18'b000011111110100001;
		14'b11101010111001:	sigmoid_prime = 18'b000011111110111100;
		14'b11101010111010:	sigmoid_prime = 18'b000011111111011000;
		14'b11101010111011:	sigmoid_prime = 18'b000011111111110011;
		14'b11101010111100:	sigmoid_prime = 18'b000100000000001111;
		14'b11101010111101:	sigmoid_prime = 18'b000100000000101011;
		14'b11101010111110:	sigmoid_prime = 18'b000100000001000111;
		14'b11101010111111:	sigmoid_prime = 18'b000100000001100011;
		14'b11101011000000:	sigmoid_prime = 18'b000100000001111110;
		14'b11101011000001:	sigmoid_prime = 18'b000100000010011010;
		14'b11101011000010:	sigmoid_prime = 18'b000100000010110110;
		14'b11101011000011:	sigmoid_prime = 18'b000100000011010010;
		14'b11101011000100:	sigmoid_prime = 18'b000100000011101110;
		14'b11101011000101:	sigmoid_prime = 18'b000100000100001010;
		14'b11101011000110:	sigmoid_prime = 18'b000100000100100110;
		14'b11101011000111:	sigmoid_prime = 18'b000100000101000011;
		14'b11101011001000:	sigmoid_prime = 18'b000100000101011111;
		14'b11101011001001:	sigmoid_prime = 18'b000100000101111011;
		14'b11101011001010:	sigmoid_prime = 18'b000100000110010111;
		14'b11101011001011:	sigmoid_prime = 18'b000100000110110100;
		14'b11101011001100:	sigmoid_prime = 18'b000100000111010000;
		14'b11101011001101:	sigmoid_prime = 18'b000100000111101100;
		14'b11101011001110:	sigmoid_prime = 18'b000100001000001001;
		14'b11101011001111:	sigmoid_prime = 18'b000100001000100101;
		14'b11101011010000:	sigmoid_prime = 18'b000100001001000010;
		14'b11101011010001:	sigmoid_prime = 18'b000100001001011110;
		14'b11101011010010:	sigmoid_prime = 18'b000100001001111011;
		14'b11101011010011:	sigmoid_prime = 18'b000100001010010111;
		14'b11101011010100:	sigmoid_prime = 18'b000100001010110100;
		14'b11101011010101:	sigmoid_prime = 18'b000100001011010001;
		14'b11101011010110:	sigmoid_prime = 18'b000100001011101110;
		14'b11101011010111:	sigmoid_prime = 18'b000100001100001010;
		14'b11101011011000:	sigmoid_prime = 18'b000100001100100111;
		14'b11101011011001:	sigmoid_prime = 18'b000100001101000100;
		14'b11101011011010:	sigmoid_prime = 18'b000100001101100001;
		14'b11101011011011:	sigmoid_prime = 18'b000100001101111110;
		14'b11101011011100:	sigmoid_prime = 18'b000100001110011011;
		14'b11101011011101:	sigmoid_prime = 18'b000100001110111000;
		14'b11101011011110:	sigmoid_prime = 18'b000100001111010101;
		14'b11101011011111:	sigmoid_prime = 18'b000100001111110010;
		14'b11101011100000:	sigmoid_prime = 18'b000100010000001111;
		14'b11101011100001:	sigmoid_prime = 18'b000100010000101100;
		14'b11101011100010:	sigmoid_prime = 18'b000100010001001010;
		14'b11101011100011:	sigmoid_prime = 18'b000100010001100111;
		14'b11101011100100:	sigmoid_prime = 18'b000100010010000100;
		14'b11101011100101:	sigmoid_prime = 18'b000100010010100001;
		14'b11101011100110:	sigmoid_prime = 18'b000100010010111111;
		14'b11101011100111:	sigmoid_prime = 18'b000100010011011100;
		14'b11101011101000:	sigmoid_prime = 18'b000100010011111010;
		14'b11101011101001:	sigmoid_prime = 18'b000100010100010111;
		14'b11101011101010:	sigmoid_prime = 18'b000100010100110101;
		14'b11101011101011:	sigmoid_prime = 18'b000100010101010010;
		14'b11101011101100:	sigmoid_prime = 18'b000100010101110000;
		14'b11101011101101:	sigmoid_prime = 18'b000100010110001110;
		14'b11101011101110:	sigmoid_prime = 18'b000100010110101011;
		14'b11101011101111:	sigmoid_prime = 18'b000100010111001001;
		14'b11101011110000:	sigmoid_prime = 18'b000100010111100111;
		14'b11101011110001:	sigmoid_prime = 18'b000100011000000101;
		14'b11101011110010:	sigmoid_prime = 18'b000100011000100010;
		14'b11101011110011:	sigmoid_prime = 18'b000100011001000000;
		14'b11101011110100:	sigmoid_prime = 18'b000100011001011110;
		14'b11101011110101:	sigmoid_prime = 18'b000100011001111100;
		14'b11101011110110:	sigmoid_prime = 18'b000100011010011010;
		14'b11101011110111:	sigmoid_prime = 18'b000100011010111000;
		14'b11101011111000:	sigmoid_prime = 18'b000100011011010110;
		14'b11101011111001:	sigmoid_prime = 18'b000100011011110101;
		14'b11101011111010:	sigmoid_prime = 18'b000100011100010011;
		14'b11101011111011:	sigmoid_prime = 18'b000100011100110001;
		14'b11101011111100:	sigmoid_prime = 18'b000100011101001111;
		14'b11101011111101:	sigmoid_prime = 18'b000100011101101110;
		14'b11101011111110:	sigmoid_prime = 18'b000100011110001100;
		14'b11101011111111:	sigmoid_prime = 18'b000100011110101010;
		14'b11101100000000:	sigmoid_prime = 18'b000100011111001001;
		14'b11101100000001:	sigmoid_prime = 18'b000100011111100111;
		14'b11101100000010:	sigmoid_prime = 18'b000100100000000110;
		14'b11101100000011:	sigmoid_prime = 18'b000100100000100100;
		14'b11101100000100:	sigmoid_prime = 18'b000100100001000011;
		14'b11101100000101:	sigmoid_prime = 18'b000100100001100010;
		14'b11101100000110:	sigmoid_prime = 18'b000100100010000000;
		14'b11101100000111:	sigmoid_prime = 18'b000100100010011111;
		14'b11101100001000:	sigmoid_prime = 18'b000100100010111110;
		14'b11101100001001:	sigmoid_prime = 18'b000100100011011100;
		14'b11101100001010:	sigmoid_prime = 18'b000100100011111011;
		14'b11101100001011:	sigmoid_prime = 18'b000100100100011010;
		14'b11101100001100:	sigmoid_prime = 18'b000100100100111001;
		14'b11101100001101:	sigmoid_prime = 18'b000100100101011000;
		14'b11101100001110:	sigmoid_prime = 18'b000100100101110111;
		14'b11101100001111:	sigmoid_prime = 18'b000100100110010110;
		14'b11101100010000:	sigmoid_prime = 18'b000100100110110101;
		14'b11101100010001:	sigmoid_prime = 18'b000100100111010100;
		14'b11101100010010:	sigmoid_prime = 18'b000100100111110011;
		14'b11101100010011:	sigmoid_prime = 18'b000100101000010011;
		14'b11101100010100:	sigmoid_prime = 18'b000100101000110010;
		14'b11101100010101:	sigmoid_prime = 18'b000100101001010001;
		14'b11101100010110:	sigmoid_prime = 18'b000100101001110000;
		14'b11101100010111:	sigmoid_prime = 18'b000100101010010000;
		14'b11101100011000:	sigmoid_prime = 18'b000100101010101111;
		14'b11101100011001:	sigmoid_prime = 18'b000100101011001111;
		14'b11101100011010:	sigmoid_prime = 18'b000100101011101110;
		14'b11101100011011:	sigmoid_prime = 18'b000100101100001110;
		14'b11101100011100:	sigmoid_prime = 18'b000100101100101101;
		14'b11101100011101:	sigmoid_prime = 18'b000100101101001101;
		14'b11101100011110:	sigmoid_prime = 18'b000100101101101101;
		14'b11101100011111:	sigmoid_prime = 18'b000100101110001100;
		14'b11101100100000:	sigmoid_prime = 18'b000100101110101100;
		14'b11101100100001:	sigmoid_prime = 18'b000100101111001100;
		14'b11101100100010:	sigmoid_prime = 18'b000100101111101100;
		14'b11101100100011:	sigmoid_prime = 18'b000100110000001011;
		14'b11101100100100:	sigmoid_prime = 18'b000100110000101011;
		14'b11101100100101:	sigmoid_prime = 18'b000100110001001011;
		14'b11101100100110:	sigmoid_prime = 18'b000100110001101011;
		14'b11101100100111:	sigmoid_prime = 18'b000100110010001011;
		14'b11101100101000:	sigmoid_prime = 18'b000100110010101011;
		14'b11101100101001:	sigmoid_prime = 18'b000100110011001011;
		14'b11101100101010:	sigmoid_prime = 18'b000100110011101100;
		14'b11101100101011:	sigmoid_prime = 18'b000100110100001100;
		14'b11101100101100:	sigmoid_prime = 18'b000100110100101100;
		14'b11101100101101:	sigmoid_prime = 18'b000100110101001100;
		14'b11101100101110:	sigmoid_prime = 18'b000100110101101101;
		14'b11101100101111:	sigmoid_prime = 18'b000100110110001101;
		14'b11101100110000:	sigmoid_prime = 18'b000100110110101101;
		14'b11101100110001:	sigmoid_prime = 18'b000100110111001110;
		14'b11101100110010:	sigmoid_prime = 18'b000100110111101110;
		14'b11101100110011:	sigmoid_prime = 18'b000100111000001111;
		14'b11101100110100:	sigmoid_prime = 18'b000100111000101111;
		14'b11101100110101:	sigmoid_prime = 18'b000100111001010000;
		14'b11101100110110:	sigmoid_prime = 18'b000100111001110001;
		14'b11101100110111:	sigmoid_prime = 18'b000100111010010001;
		14'b11101100111000:	sigmoid_prime = 18'b000100111010110010;
		14'b11101100111001:	sigmoid_prime = 18'b000100111011010011;
		14'b11101100111010:	sigmoid_prime = 18'b000100111011110100;
		14'b11101100111011:	sigmoid_prime = 18'b000100111100010100;
		14'b11101100111100:	sigmoid_prime = 18'b000100111100110101;
		14'b11101100111101:	sigmoid_prime = 18'b000100111101010110;
		14'b11101100111110:	sigmoid_prime = 18'b000100111101110111;
		14'b11101100111111:	sigmoid_prime = 18'b000100111110011000;
		14'b11101101000000:	sigmoid_prime = 18'b000100111110111001;
		14'b11101101000001:	sigmoid_prime = 18'b000100111111011010;
		14'b11101101000010:	sigmoid_prime = 18'b000100111111111100;
		14'b11101101000011:	sigmoid_prime = 18'b000101000000011101;
		14'b11101101000100:	sigmoid_prime = 18'b000101000000111110;
		14'b11101101000101:	sigmoid_prime = 18'b000101000001011111;
		14'b11101101000110:	sigmoid_prime = 18'b000101000010000001;
		14'b11101101000111:	sigmoid_prime = 18'b000101000010100010;
		14'b11101101001000:	sigmoid_prime = 18'b000101000011000011;
		14'b11101101001001:	sigmoid_prime = 18'b000101000011100101;
		14'b11101101001010:	sigmoid_prime = 18'b000101000100000110;
		14'b11101101001011:	sigmoid_prime = 18'b000101000100101000;
		14'b11101101001100:	sigmoid_prime = 18'b000101000101001001;
		14'b11101101001101:	sigmoid_prime = 18'b000101000101101011;
		14'b11101101001110:	sigmoid_prime = 18'b000101000110001100;
		14'b11101101001111:	sigmoid_prime = 18'b000101000110101110;
		14'b11101101010000:	sigmoid_prime = 18'b000101000111010000;
		14'b11101101010001:	sigmoid_prime = 18'b000101000111110010;
		14'b11101101010010:	sigmoid_prime = 18'b000101001000010011;
		14'b11101101010011:	sigmoid_prime = 18'b000101001000110101;
		14'b11101101010100:	sigmoid_prime = 18'b000101001001010111;
		14'b11101101010101:	sigmoid_prime = 18'b000101001001111001;
		14'b11101101010110:	sigmoid_prime = 18'b000101001010011011;
		14'b11101101010111:	sigmoid_prime = 18'b000101001010111101;
		14'b11101101011000:	sigmoid_prime = 18'b000101001011011111;
		14'b11101101011001:	sigmoid_prime = 18'b000101001100000001;
		14'b11101101011010:	sigmoid_prime = 18'b000101001100100011;
		14'b11101101011011:	sigmoid_prime = 18'b000101001101000110;
		14'b11101101011100:	sigmoid_prime = 18'b000101001101101000;
		14'b11101101011101:	sigmoid_prime = 18'b000101001110001010;
		14'b11101101011110:	sigmoid_prime = 18'b000101001110101100;
		14'b11101101011111:	sigmoid_prime = 18'b000101001111001111;
		14'b11101101100000:	sigmoid_prime = 18'b000101001111110001;
		14'b11101101100001:	sigmoid_prime = 18'b000101010000010100;
		14'b11101101100010:	sigmoid_prime = 18'b000101010000110110;
		14'b11101101100011:	sigmoid_prime = 18'b000101010001011000;
		14'b11101101100100:	sigmoid_prime = 18'b000101010001111011;
		14'b11101101100101:	sigmoid_prime = 18'b000101010010011110;
		14'b11101101100110:	sigmoid_prime = 18'b000101010011000000;
		14'b11101101100111:	sigmoid_prime = 18'b000101010011100011;
		14'b11101101101000:	sigmoid_prime = 18'b000101010100000110;
		14'b11101101101001:	sigmoid_prime = 18'b000101010100101000;
		14'b11101101101010:	sigmoid_prime = 18'b000101010101001011;
		14'b11101101101011:	sigmoid_prime = 18'b000101010101101110;
		14'b11101101101100:	sigmoid_prime = 18'b000101010110010001;
		14'b11101101101101:	sigmoid_prime = 18'b000101010110110100;
		14'b11101101101110:	sigmoid_prime = 18'b000101010111010111;
		14'b11101101101111:	sigmoid_prime = 18'b000101010111111010;
		14'b11101101110000:	sigmoid_prime = 18'b000101011000011101;
		14'b11101101110001:	sigmoid_prime = 18'b000101011001000000;
		14'b11101101110010:	sigmoid_prime = 18'b000101011001100011;
		14'b11101101110011:	sigmoid_prime = 18'b000101011010000110;
		14'b11101101110100:	sigmoid_prime = 18'b000101011010101010;
		14'b11101101110101:	sigmoid_prime = 18'b000101011011001101;
		14'b11101101110110:	sigmoid_prime = 18'b000101011011110000;
		14'b11101101110111:	sigmoid_prime = 18'b000101011100010100;
		14'b11101101111000:	sigmoid_prime = 18'b000101011100110111;
		14'b11101101111001:	sigmoid_prime = 18'b000101011101011010;
		14'b11101101111010:	sigmoid_prime = 18'b000101011101111110;
		14'b11101101111011:	sigmoid_prime = 18'b000101011110100001;
		14'b11101101111100:	sigmoid_prime = 18'b000101011111000101;
		14'b11101101111101:	sigmoid_prime = 18'b000101011111101000;
		14'b11101101111110:	sigmoid_prime = 18'b000101100000001100;
		14'b11101101111111:	sigmoid_prime = 18'b000101100000110000;
		14'b11101110000000:	sigmoid_prime = 18'b000101100001010100;
		14'b11101110000001:	sigmoid_prime = 18'b000101100001110111;
		14'b11101110000010:	sigmoid_prime = 18'b000101100010011011;
		14'b11101110000011:	sigmoid_prime = 18'b000101100010111111;
		14'b11101110000100:	sigmoid_prime = 18'b000101100011100011;
		14'b11101110000101:	sigmoid_prime = 18'b000101100100000111;
		14'b11101110000110:	sigmoid_prime = 18'b000101100100101011;
		14'b11101110000111:	sigmoid_prime = 18'b000101100101001111;
		14'b11101110001000:	sigmoid_prime = 18'b000101100101110011;
		14'b11101110001001:	sigmoid_prime = 18'b000101100110010111;
		14'b11101110001010:	sigmoid_prime = 18'b000101100110111011;
		14'b11101110001011:	sigmoid_prime = 18'b000101100111011111;
		14'b11101110001100:	sigmoid_prime = 18'b000101101000000011;
		14'b11101110001101:	sigmoid_prime = 18'b000101101000101000;
		14'b11101110001110:	sigmoid_prime = 18'b000101101001001100;
		14'b11101110001111:	sigmoid_prime = 18'b000101101001110000;
		14'b11101110010000:	sigmoid_prime = 18'b000101101010010101;
		14'b11101110010001:	sigmoid_prime = 18'b000101101010111001;
		14'b11101110010010:	sigmoid_prime = 18'b000101101011011110;
		14'b11101110010011:	sigmoid_prime = 18'b000101101100000010;
		14'b11101110010100:	sigmoid_prime = 18'b000101101100100111;
		14'b11101110010101:	sigmoid_prime = 18'b000101101101001011;
		14'b11101110010110:	sigmoid_prime = 18'b000101101101110000;
		14'b11101110010111:	sigmoid_prime = 18'b000101101110010101;
		14'b11101110011000:	sigmoid_prime = 18'b000101101110111001;
		14'b11101110011001:	sigmoid_prime = 18'b000101101111011110;
		14'b11101110011010:	sigmoid_prime = 18'b000101110000000011;
		14'b11101110011011:	sigmoid_prime = 18'b000101110000101000;
		14'b11101110011100:	sigmoid_prime = 18'b000101110001001101;
		14'b11101110011101:	sigmoid_prime = 18'b000101110001110001;
		14'b11101110011110:	sigmoid_prime = 18'b000101110010010110;
		14'b11101110011111:	sigmoid_prime = 18'b000101110010111011;
		14'b11101110100000:	sigmoid_prime = 18'b000101110011100001;
		14'b11101110100001:	sigmoid_prime = 18'b000101110100000110;
		14'b11101110100010:	sigmoid_prime = 18'b000101110100101011;
		14'b11101110100011:	sigmoid_prime = 18'b000101110101010000;
		14'b11101110100100:	sigmoid_prime = 18'b000101110101110101;
		14'b11101110100101:	sigmoid_prime = 18'b000101110110011010;
		14'b11101110100110:	sigmoid_prime = 18'b000101110111000000;
		14'b11101110100111:	sigmoid_prime = 18'b000101110111100101;
		14'b11101110101000:	sigmoid_prime = 18'b000101111000001010;
		14'b11101110101001:	sigmoid_prime = 18'b000101111000110000;
		14'b11101110101010:	sigmoid_prime = 18'b000101111001010101;
		14'b11101110101011:	sigmoid_prime = 18'b000101111001111011;
		14'b11101110101100:	sigmoid_prime = 18'b000101111010100000;
		14'b11101110101101:	sigmoid_prime = 18'b000101111011000110;
		14'b11101110101110:	sigmoid_prime = 18'b000101111011101100;
		14'b11101110101111:	sigmoid_prime = 18'b000101111100010001;
		14'b11101110110000:	sigmoid_prime = 18'b000101111100110111;
		14'b11101110110001:	sigmoid_prime = 18'b000101111101011101;
		14'b11101110110010:	sigmoid_prime = 18'b000101111110000010;
		14'b11101110110011:	sigmoid_prime = 18'b000101111110101000;
		14'b11101110110100:	sigmoid_prime = 18'b000101111111001110;
		14'b11101110110101:	sigmoid_prime = 18'b000101111111110100;
		14'b11101110110110:	sigmoid_prime = 18'b000110000000011010;
		14'b11101110110111:	sigmoid_prime = 18'b000110000001000000;
		14'b11101110111000:	sigmoid_prime = 18'b000110000001100110;
		14'b11101110111001:	sigmoid_prime = 18'b000110000010001100;
		14'b11101110111010:	sigmoid_prime = 18'b000110000010110010;
		14'b11101110111011:	sigmoid_prime = 18'b000110000011011000;
		14'b11101110111100:	sigmoid_prime = 18'b000110000011111111;
		14'b11101110111101:	sigmoid_prime = 18'b000110000100100101;
		14'b11101110111110:	sigmoid_prime = 18'b000110000101001011;
		14'b11101110111111:	sigmoid_prime = 18'b000110000101110001;
		14'b11101111000000:	sigmoid_prime = 18'b000110000110011000;
		14'b11101111000001:	sigmoid_prime = 18'b000110000110111110;
		14'b11101111000010:	sigmoid_prime = 18'b000110000111100101;
		14'b11101111000011:	sigmoid_prime = 18'b000110001000001011;
		14'b11101111000100:	sigmoid_prime = 18'b000110001000110010;
		14'b11101111000101:	sigmoid_prime = 18'b000110001001011000;
		14'b11101111000110:	sigmoid_prime = 18'b000110001001111111;
		14'b11101111000111:	sigmoid_prime = 18'b000110001010100110;
		14'b11101111001000:	sigmoid_prime = 18'b000110001011001100;
		14'b11101111001001:	sigmoid_prime = 18'b000110001011110011;
		14'b11101111001010:	sigmoid_prime = 18'b000110001100011010;
		14'b11101111001011:	sigmoid_prime = 18'b000110001101000001;
		14'b11101111001100:	sigmoid_prime = 18'b000110001101100111;
		14'b11101111001101:	sigmoid_prime = 18'b000110001110001110;
		14'b11101111001110:	sigmoid_prime = 18'b000110001110110101;
		14'b11101111001111:	sigmoid_prime = 18'b000110001111011100;
		14'b11101111010000:	sigmoid_prime = 18'b000110010000000011;
		14'b11101111010001:	sigmoid_prime = 18'b000110010000101010;
		14'b11101111010010:	sigmoid_prime = 18'b000110010001010001;
		14'b11101111010011:	sigmoid_prime = 18'b000110010001111001;
		14'b11101111010100:	sigmoid_prime = 18'b000110010010100000;
		14'b11101111010101:	sigmoid_prime = 18'b000110010011000111;
		14'b11101111010110:	sigmoid_prime = 18'b000110010011101110;
		14'b11101111010111:	sigmoid_prime = 18'b000110010100010101;
		14'b11101111011000:	sigmoid_prime = 18'b000110010100111101;
		14'b11101111011001:	sigmoid_prime = 18'b000110010101100100;
		14'b11101111011010:	sigmoid_prime = 18'b000110010110001100;
		14'b11101111011011:	sigmoid_prime = 18'b000110010110110011;
		14'b11101111011100:	sigmoid_prime = 18'b000110010111011011;
		14'b11101111011101:	sigmoid_prime = 18'b000110011000000010;
		14'b11101111011110:	sigmoid_prime = 18'b000110011000101010;
		14'b11101111011111:	sigmoid_prime = 18'b000110011001010001;
		14'b11101111100000:	sigmoid_prime = 18'b000110011001111001;
		14'b11101111100001:	sigmoid_prime = 18'b000110011010100001;
		14'b11101111100010:	sigmoid_prime = 18'b000110011011001000;
		14'b11101111100011:	sigmoid_prime = 18'b000110011011110000;
		14'b11101111100100:	sigmoid_prime = 18'b000110011100011000;
		14'b11101111100101:	sigmoid_prime = 18'b000110011101000000;
		14'b11101111100110:	sigmoid_prime = 18'b000110011101101000;
		14'b11101111100111:	sigmoid_prime = 18'b000110011110010000;
		14'b11101111101000:	sigmoid_prime = 18'b000110011110111000;
		14'b11101111101001:	sigmoid_prime = 18'b000110011111100000;
		14'b11101111101010:	sigmoid_prime = 18'b000110100000001000;
		14'b11101111101011:	sigmoid_prime = 18'b000110100000110000;
		14'b11101111101100:	sigmoid_prime = 18'b000110100001011000;
		14'b11101111101101:	sigmoid_prime = 18'b000110100010000000;
		14'b11101111101110:	sigmoid_prime = 18'b000110100010101000;
		14'b11101111101111:	sigmoid_prime = 18'b000110100011010001;
		14'b11101111110000:	sigmoid_prime = 18'b000110100011111001;
		14'b11101111110001:	sigmoid_prime = 18'b000110100100100001;
		14'b11101111110010:	sigmoid_prime = 18'b000110100101001010;
		14'b11101111110011:	sigmoid_prime = 18'b000110100101110010;
		14'b11101111110100:	sigmoid_prime = 18'b000110100110011010;
		14'b11101111110101:	sigmoid_prime = 18'b000110100111000011;
		14'b11101111110110:	sigmoid_prime = 18'b000110100111101011;
		14'b11101111110111:	sigmoid_prime = 18'b000110101000010100;
		14'b11101111111000:	sigmoid_prime = 18'b000110101000111101;
		14'b11101111111001:	sigmoid_prime = 18'b000110101001100101;
		14'b11101111111010:	sigmoid_prime = 18'b000110101010001110;
		14'b11101111111011:	sigmoid_prime = 18'b000110101010110111;
		14'b11101111111100:	sigmoid_prime = 18'b000110101011011111;
		14'b11101111111101:	sigmoid_prime = 18'b000110101100001000;
		14'b11101111111110:	sigmoid_prime = 18'b000110101100110001;
		14'b11101111111111:	sigmoid_prime = 18'b000110101101011010;
		14'b11110000000000:	sigmoid_prime = 18'b000110101110000011;
		14'b11110000000001:	sigmoid_prime = 18'b000110101110101100;
		14'b11110000000010:	sigmoid_prime = 18'b000110101111010101;
		14'b11110000000011:	sigmoid_prime = 18'b000110101111111110;
		14'b11110000000100:	sigmoid_prime = 18'b000110110000100111;
		14'b11110000000101:	sigmoid_prime = 18'b000110110001010000;
		14'b11110000000110:	sigmoid_prime = 18'b000110110001111001;
		14'b11110000000111:	sigmoid_prime = 18'b000110110010100010;
		14'b11110000001000:	sigmoid_prime = 18'b000110110011001100;
		14'b11110000001001:	sigmoid_prime = 18'b000110110011110101;
		14'b11110000001010:	sigmoid_prime = 18'b000110110100011110;
		14'b11110000001011:	sigmoid_prime = 18'b000110110101001000;
		14'b11110000001100:	sigmoid_prime = 18'b000110110101110001;
		14'b11110000001101:	sigmoid_prime = 18'b000110110110011010;
		14'b11110000001110:	sigmoid_prime = 18'b000110110111000100;
		14'b11110000001111:	sigmoid_prime = 18'b000110110111101101;
		14'b11110000010000:	sigmoid_prime = 18'b000110111000010111;
		14'b11110000010001:	sigmoid_prime = 18'b000110111001000001;
		14'b11110000010010:	sigmoid_prime = 18'b000110111001101010;
		14'b11110000010011:	sigmoid_prime = 18'b000110111010010100;
		14'b11110000010100:	sigmoid_prime = 18'b000110111010111101;
		14'b11110000010101:	sigmoid_prime = 18'b000110111011100111;
		14'b11110000010110:	sigmoid_prime = 18'b000110111100010001;
		14'b11110000010111:	sigmoid_prime = 18'b000110111100111011;
		14'b11110000011000:	sigmoid_prime = 18'b000110111101100101;
		14'b11110000011001:	sigmoid_prime = 18'b000110111110001110;
		14'b11110000011010:	sigmoid_prime = 18'b000110111110111000;
		14'b11110000011011:	sigmoid_prime = 18'b000110111111100010;
		14'b11110000011100:	sigmoid_prime = 18'b000111000000001100;
		14'b11110000011101:	sigmoid_prime = 18'b000111000000110110;
		14'b11110000011110:	sigmoid_prime = 18'b000111000001100000;
		14'b11110000011111:	sigmoid_prime = 18'b000111000010001011;
		14'b11110000100000:	sigmoid_prime = 18'b000111000010110101;
		14'b11110000100001:	sigmoid_prime = 18'b000111000011011111;
		14'b11110000100010:	sigmoid_prime = 18'b000111000100001001;
		14'b11110000100011:	sigmoid_prime = 18'b000111000100110011;
		14'b11110000100100:	sigmoid_prime = 18'b000111000101011110;
		14'b11110000100101:	sigmoid_prime = 18'b000111000110001000;
		14'b11110000100110:	sigmoid_prime = 18'b000111000110110010;
		14'b11110000100111:	sigmoid_prime = 18'b000111000111011101;
		14'b11110000101000:	sigmoid_prime = 18'b000111001000000111;
		14'b11110000101001:	sigmoid_prime = 18'b000111001000110010;
		14'b11110000101010:	sigmoid_prime = 18'b000111001001011100;
		14'b11110000101011:	sigmoid_prime = 18'b000111001010000111;
		14'b11110000101100:	sigmoid_prime = 18'b000111001010110001;
		14'b11110000101101:	sigmoid_prime = 18'b000111001011011100;
		14'b11110000101110:	sigmoid_prime = 18'b000111001100000111;
		14'b11110000101111:	sigmoid_prime = 18'b000111001100110001;
		14'b11110000110000:	sigmoid_prime = 18'b000111001101011100;
		14'b11110000110001:	sigmoid_prime = 18'b000111001110000111;
		14'b11110000110010:	sigmoid_prime = 18'b000111001110110010;
		14'b11110000110011:	sigmoid_prime = 18'b000111001111011100;
		14'b11110000110100:	sigmoid_prime = 18'b000111010000000111;
		14'b11110000110101:	sigmoid_prime = 18'b000111010000110010;
		14'b11110000110110:	sigmoid_prime = 18'b000111010001011101;
		14'b11110000110111:	sigmoid_prime = 18'b000111010010001000;
		14'b11110000111000:	sigmoid_prime = 18'b000111010010110011;
		14'b11110000111001:	sigmoid_prime = 18'b000111010011011110;
		14'b11110000111010:	sigmoid_prime = 18'b000111010100001001;
		14'b11110000111011:	sigmoid_prime = 18'b000111010100110101;
		14'b11110000111100:	sigmoid_prime = 18'b000111010101100000;
		14'b11110000111101:	sigmoid_prime = 18'b000111010110001011;
		14'b11110000111110:	sigmoid_prime = 18'b000111010110110110;
		14'b11110000111111:	sigmoid_prime = 18'b000111010111100001;
		14'b11110001000000:	sigmoid_prime = 18'b000111011000001101;
		14'b11110001000001:	sigmoid_prime = 18'b000111011000111000;
		14'b11110001000010:	sigmoid_prime = 18'b000111011001100011;
		14'b11110001000011:	sigmoid_prime = 18'b000111011010001111;
		14'b11110001000100:	sigmoid_prime = 18'b000111011010111010;
		14'b11110001000101:	sigmoid_prime = 18'b000111011011100110;
		14'b11110001000110:	sigmoid_prime = 18'b000111011100010001;
		14'b11110001000111:	sigmoid_prime = 18'b000111011100111101;
		14'b11110001001000:	sigmoid_prime = 18'b000111011101101000;
		14'b11110001001001:	sigmoid_prime = 18'b000111011110010100;
		14'b11110001001010:	sigmoid_prime = 18'b000111011111000000;
		14'b11110001001011:	sigmoid_prime = 18'b000111011111101011;
		14'b11110001001100:	sigmoid_prime = 18'b000111100000010111;
		14'b11110001001101:	sigmoid_prime = 18'b000111100001000011;
		14'b11110001001110:	sigmoid_prime = 18'b000111100001101111;
		14'b11110001001111:	sigmoid_prime = 18'b000111100010011011;
		14'b11110001010000:	sigmoid_prime = 18'b000111100011000110;
		14'b11110001010001:	sigmoid_prime = 18'b000111100011110010;
		14'b11110001010010:	sigmoid_prime = 18'b000111100100011110;
		14'b11110001010011:	sigmoid_prime = 18'b000111100101001010;
		14'b11110001010100:	sigmoid_prime = 18'b000111100101110110;
		14'b11110001010101:	sigmoid_prime = 18'b000111100110100010;
		14'b11110001010110:	sigmoid_prime = 18'b000111100111001110;
		14'b11110001010111:	sigmoid_prime = 18'b000111100111111011;
		14'b11110001011000:	sigmoid_prime = 18'b000111101000100111;
		14'b11110001011001:	sigmoid_prime = 18'b000111101001010011;
		14'b11110001011010:	sigmoid_prime = 18'b000111101001111111;
		14'b11110001011011:	sigmoid_prime = 18'b000111101010101011;
		14'b11110001011100:	sigmoid_prime = 18'b000111101011011000;
		14'b11110001011101:	sigmoid_prime = 18'b000111101100000100;
		14'b11110001011110:	sigmoid_prime = 18'b000111101100110000;
		14'b11110001011111:	sigmoid_prime = 18'b000111101101011101;
		14'b11110001100000:	sigmoid_prime = 18'b000111101110001001;
		14'b11110001100001:	sigmoid_prime = 18'b000111101110110110;
		14'b11110001100010:	sigmoid_prime = 18'b000111101111100010;
		14'b11110001100011:	sigmoid_prime = 18'b000111110000001111;
		14'b11110001100100:	sigmoid_prime = 18'b000111110000111011;
		14'b11110001100101:	sigmoid_prime = 18'b000111110001101000;
		14'b11110001100110:	sigmoid_prime = 18'b000111110010010100;
		14'b11110001100111:	sigmoid_prime = 18'b000111110011000001;
		14'b11110001101000:	sigmoid_prime = 18'b000111110011101110;
		14'b11110001101001:	sigmoid_prime = 18'b000111110100011010;
		14'b11110001101010:	sigmoid_prime = 18'b000111110101000111;
		14'b11110001101011:	sigmoid_prime = 18'b000111110101110100;
		14'b11110001101100:	sigmoid_prime = 18'b000111110110100001;
		14'b11110001101101:	sigmoid_prime = 18'b000111110111001101;
		14'b11110001101110:	sigmoid_prime = 18'b000111110111111010;
		14'b11110001101111:	sigmoid_prime = 18'b000111111000100111;
		14'b11110001110000:	sigmoid_prime = 18'b000111111001010100;
		14'b11110001110001:	sigmoid_prime = 18'b000111111010000001;
		14'b11110001110010:	sigmoid_prime = 18'b000111111010101110;
		14'b11110001110011:	sigmoid_prime = 18'b000111111011011011;
		14'b11110001110100:	sigmoid_prime = 18'b000111111100001000;
		14'b11110001110101:	sigmoid_prime = 18'b000111111100110101;
		14'b11110001110110:	sigmoid_prime = 18'b000111111101100010;
		14'b11110001110111:	sigmoid_prime = 18'b000111111110010000;
		14'b11110001111000:	sigmoid_prime = 18'b000111111110111101;
		14'b11110001111001:	sigmoid_prime = 18'b000111111111101010;
		14'b11110001111010:	sigmoid_prime = 18'b001000000000010111;
		14'b11110001111011:	sigmoid_prime = 18'b001000000001000101;
		14'b11110001111100:	sigmoid_prime = 18'b001000000001110010;
		14'b11110001111101:	sigmoid_prime = 18'b001000000010011111;
		14'b11110001111110:	sigmoid_prime = 18'b001000000011001101;
		14'b11110001111111:	sigmoid_prime = 18'b001000000011111010;
		14'b11110010000000:	sigmoid_prime = 18'b001000000100101000;
		14'b11110010000001:	sigmoid_prime = 18'b001000000101010101;
		14'b11110010000010:	sigmoid_prime = 18'b001000000110000010;
		14'b11110010000011:	sigmoid_prime = 18'b001000000110110000;
		14'b11110010000100:	sigmoid_prime = 18'b001000000111011110;
		14'b11110010000101:	sigmoid_prime = 18'b001000001000001011;
		14'b11110010000110:	sigmoid_prime = 18'b001000001000111001;
		14'b11110010000111:	sigmoid_prime = 18'b001000001001100110;
		14'b11110010001000:	sigmoid_prime = 18'b001000001010010100;
		14'b11110010001001:	sigmoid_prime = 18'b001000001011000010;
		14'b11110010001010:	sigmoid_prime = 18'b001000001011110000;
		14'b11110010001011:	sigmoid_prime = 18'b001000001100011101;
		14'b11110010001100:	sigmoid_prime = 18'b001000001101001011;
		14'b11110010001101:	sigmoid_prime = 18'b001000001101111001;
		14'b11110010001110:	sigmoid_prime = 18'b001000001110100111;
		14'b11110010001111:	sigmoid_prime = 18'b001000001111010101;
		14'b11110010010000:	sigmoid_prime = 18'b001000010000000011;
		14'b11110010010001:	sigmoid_prime = 18'b001000010000110001;
		14'b11110010010010:	sigmoid_prime = 18'b001000010001011111;
		14'b11110010010011:	sigmoid_prime = 18'b001000010010001101;
		14'b11110010010100:	sigmoid_prime = 18'b001000010010111011;
		14'b11110010010101:	sigmoid_prime = 18'b001000010011101001;
		14'b11110010010110:	sigmoid_prime = 18'b001000010100010111;
		14'b11110010010111:	sigmoid_prime = 18'b001000010101000101;
		14'b11110010011000:	sigmoid_prime = 18'b001000010101110011;
		14'b11110010011001:	sigmoid_prime = 18'b001000010110100001;
		14'b11110010011010:	sigmoid_prime = 18'b001000010111001111;
		14'b11110010011011:	sigmoid_prime = 18'b001000010111111110;
		14'b11110010011100:	sigmoid_prime = 18'b001000011000101100;
		14'b11110010011101:	sigmoid_prime = 18'b001000011001011010;
		14'b11110010011110:	sigmoid_prime = 18'b001000011010001001;
		14'b11110010011111:	sigmoid_prime = 18'b001000011010110111;
		14'b11110010100000:	sigmoid_prime = 18'b001000011011100101;
		14'b11110010100001:	sigmoid_prime = 18'b001000011100010100;
		14'b11110010100010:	sigmoid_prime = 18'b001000011101000010;
		14'b11110010100011:	sigmoid_prime = 18'b001000011101110001;
		14'b11110010100100:	sigmoid_prime = 18'b001000011110011111;
		14'b11110010100101:	sigmoid_prime = 18'b001000011111001110;
		14'b11110010100110:	sigmoid_prime = 18'b001000011111111100;
		14'b11110010100111:	sigmoid_prime = 18'b001000100000101011;
		14'b11110010101000:	sigmoid_prime = 18'b001000100001011001;
		14'b11110010101001:	sigmoid_prime = 18'b001000100010001000;
		14'b11110010101010:	sigmoid_prime = 18'b001000100010110111;
		14'b11110010101011:	sigmoid_prime = 18'b001000100011100101;
		14'b11110010101100:	sigmoid_prime = 18'b001000100100010100;
		14'b11110010101101:	sigmoid_prime = 18'b001000100101000011;
		14'b11110010101110:	sigmoid_prime = 18'b001000100101110001;
		14'b11110010101111:	sigmoid_prime = 18'b001000100110100000;
		14'b11110010110000:	sigmoid_prime = 18'b001000100111001111;
		14'b11110010110001:	sigmoid_prime = 18'b001000100111111110;
		14'b11110010110010:	sigmoid_prime = 18'b001000101000101101;
		14'b11110010110011:	sigmoid_prime = 18'b001000101001011100;
		14'b11110010110100:	sigmoid_prime = 18'b001000101010001011;
		14'b11110010110101:	sigmoid_prime = 18'b001000101010111001;
		14'b11110010110110:	sigmoid_prime = 18'b001000101011101000;
		14'b11110010110111:	sigmoid_prime = 18'b001000101100010111;
		14'b11110010111000:	sigmoid_prime = 18'b001000101101000110;
		14'b11110010111001:	sigmoid_prime = 18'b001000101101110101;
		14'b11110010111010:	sigmoid_prime = 18'b001000101110100101;
		14'b11110010111011:	sigmoid_prime = 18'b001000101111010100;
		14'b11110010111100:	sigmoid_prime = 18'b001000110000000011;
		14'b11110010111101:	sigmoid_prime = 18'b001000110000110010;
		14'b11110010111110:	sigmoid_prime = 18'b001000110001100001;
		14'b11110010111111:	sigmoid_prime = 18'b001000110010010000;
		14'b11110011000000:	sigmoid_prime = 18'b001000110010111111;
		14'b11110011000001:	sigmoid_prime = 18'b001000110011101111;
		14'b11110011000010:	sigmoid_prime = 18'b001000110100011110;
		14'b11110011000011:	sigmoid_prime = 18'b001000110101001101;
		14'b11110011000100:	sigmoid_prime = 18'b001000110101111100;
		14'b11110011000101:	sigmoid_prime = 18'b001000110110101100;
		14'b11110011000110:	sigmoid_prime = 18'b001000110111011011;
		14'b11110011000111:	sigmoid_prime = 18'b001000111000001011;
		14'b11110011001000:	sigmoid_prime = 18'b001000111000111010;
		14'b11110011001001:	sigmoid_prime = 18'b001000111001101001;
		14'b11110011001010:	sigmoid_prime = 18'b001000111010011001;
		14'b11110011001011:	sigmoid_prime = 18'b001000111011001000;
		14'b11110011001100:	sigmoid_prime = 18'b001000111011111000;
		14'b11110011001101:	sigmoid_prime = 18'b001000111100100111;
		14'b11110011001110:	sigmoid_prime = 18'b001000111101010111;
		14'b11110011001111:	sigmoid_prime = 18'b001000111110000110;
		14'b11110011010000:	sigmoid_prime = 18'b001000111110110110;
		14'b11110011010001:	sigmoid_prime = 18'b001000111111100110;
		14'b11110011010010:	sigmoid_prime = 18'b001001000000010101;
		14'b11110011010011:	sigmoid_prime = 18'b001001000001000101;
		14'b11110011010100:	sigmoid_prime = 18'b001001000001110100;
		14'b11110011010101:	sigmoid_prime = 18'b001001000010100100;
		14'b11110011010110:	sigmoid_prime = 18'b001001000011010100;
		14'b11110011010111:	sigmoid_prime = 18'b001001000100000100;
		14'b11110011011000:	sigmoid_prime = 18'b001001000100110011;
		14'b11110011011001:	sigmoid_prime = 18'b001001000101100011;
		14'b11110011011010:	sigmoid_prime = 18'b001001000110010011;
		14'b11110011011011:	sigmoid_prime = 18'b001001000111000011;
		14'b11110011011100:	sigmoid_prime = 18'b001001000111110011;
		14'b11110011011101:	sigmoid_prime = 18'b001001001000100010;
		14'b11110011011110:	sigmoid_prime = 18'b001001001001010010;
		14'b11110011011111:	sigmoid_prime = 18'b001001001010000010;
		14'b11110011100000:	sigmoid_prime = 18'b001001001010110010;
		14'b11110011100001:	sigmoid_prime = 18'b001001001011100010;
		14'b11110011100010:	sigmoid_prime = 18'b001001001100010010;
		14'b11110011100011:	sigmoid_prime = 18'b001001001101000010;
		14'b11110011100100:	sigmoid_prime = 18'b001001001101110010;
		14'b11110011100101:	sigmoid_prime = 18'b001001001110100010;
		14'b11110011100110:	sigmoid_prime = 18'b001001001111010010;
		14'b11110011100111:	sigmoid_prime = 18'b001001010000000010;
		14'b11110011101000:	sigmoid_prime = 18'b001001010000110010;
		14'b11110011101001:	sigmoid_prime = 18'b001001010001100010;
		14'b11110011101010:	sigmoid_prime = 18'b001001010010010010;
		14'b11110011101011:	sigmoid_prime = 18'b001001010011000010;
		14'b11110011101100:	sigmoid_prime = 18'b001001010011110011;
		14'b11110011101101:	sigmoid_prime = 18'b001001010100100011;
		14'b11110011101110:	sigmoid_prime = 18'b001001010101010011;
		14'b11110011101111:	sigmoid_prime = 18'b001001010110000011;
		14'b11110011110000:	sigmoid_prime = 18'b001001010110110011;
		14'b11110011110001:	sigmoid_prime = 18'b001001010111100100;
		14'b11110011110010:	sigmoid_prime = 18'b001001011000010100;
		14'b11110011110011:	sigmoid_prime = 18'b001001011001000100;
		14'b11110011110100:	sigmoid_prime = 18'b001001011001110100;
		14'b11110011110101:	sigmoid_prime = 18'b001001011010100101;
		14'b11110011110110:	sigmoid_prime = 18'b001001011011010101;
		14'b11110011110111:	sigmoid_prime = 18'b001001011100000101;
		14'b11110011111000:	sigmoid_prime = 18'b001001011100110110;
		14'b11110011111001:	sigmoid_prime = 18'b001001011101100110;
		14'b11110011111010:	sigmoid_prime = 18'b001001011110010111;
		14'b11110011111011:	sigmoid_prime = 18'b001001011111000111;
		14'b11110011111100:	sigmoid_prime = 18'b001001011111110111;
		14'b11110011111101:	sigmoid_prime = 18'b001001100000101000;
		14'b11110011111110:	sigmoid_prime = 18'b001001100001011000;
		14'b11110011111111:	sigmoid_prime = 18'b001001100010001001;
		14'b11110100000000:	sigmoid_prime = 18'b001001100010111001;
		14'b11110100000001:	sigmoid_prime = 18'b001001100011101010;
		14'b11110100000010:	sigmoid_prime = 18'b001001100100011010;
		14'b11110100000011:	sigmoid_prime = 18'b001001100101001011;
		14'b11110100000100:	sigmoid_prime = 18'b001001100101111011;
		14'b11110100000101:	sigmoid_prime = 18'b001001100110101100;
		14'b11110100000110:	sigmoid_prime = 18'b001001100111011101;
		14'b11110100000111:	sigmoid_prime = 18'b001001101000001101;
		14'b11110100001000:	sigmoid_prime = 18'b001001101000111110;
		14'b11110100001001:	sigmoid_prime = 18'b001001101001101110;
		14'b11110100001010:	sigmoid_prime = 18'b001001101010011111;
		14'b11110100001011:	sigmoid_prime = 18'b001001101011010000;
		14'b11110100001100:	sigmoid_prime = 18'b001001101100000000;
		14'b11110100001101:	sigmoid_prime = 18'b001001101100110001;
		14'b11110100001110:	sigmoid_prime = 18'b001001101101100010;
		14'b11110100001111:	sigmoid_prime = 18'b001001101110010011;
		14'b11110100010000:	sigmoid_prime = 18'b001001101111000011;
		14'b11110100010001:	sigmoid_prime = 18'b001001101111110100;
		14'b11110100010010:	sigmoid_prime = 18'b001001110000100101;
		14'b11110100010011:	sigmoid_prime = 18'b001001110001010110;
		14'b11110100010100:	sigmoid_prime = 18'b001001110010000110;
		14'b11110100010101:	sigmoid_prime = 18'b001001110010110111;
		14'b11110100010110:	sigmoid_prime = 18'b001001110011101000;
		14'b11110100010111:	sigmoid_prime = 18'b001001110100011001;
		14'b11110100011000:	sigmoid_prime = 18'b001001110101001010;
		14'b11110100011001:	sigmoid_prime = 18'b001001110101111010;
		14'b11110100011010:	sigmoid_prime = 18'b001001110110101011;
		14'b11110100011011:	sigmoid_prime = 18'b001001110111011100;
		14'b11110100011100:	sigmoid_prime = 18'b001001111000001101;
		14'b11110100011101:	sigmoid_prime = 18'b001001111000111110;
		14'b11110100011110:	sigmoid_prime = 18'b001001111001101111;
		14'b11110100011111:	sigmoid_prime = 18'b001001111010100000;
		14'b11110100100000:	sigmoid_prime = 18'b001001111011010001;
		14'b11110100100001:	sigmoid_prime = 18'b001001111100000010;
		14'b11110100100010:	sigmoid_prime = 18'b001001111100110010;
		14'b11110100100011:	sigmoid_prime = 18'b001001111101100011;
		14'b11110100100100:	sigmoid_prime = 18'b001001111110010100;
		14'b11110100100101:	sigmoid_prime = 18'b001001111111000101;
		14'b11110100100110:	sigmoid_prime = 18'b001001111111110110;
		14'b11110100100111:	sigmoid_prime = 18'b001010000000100111;
		14'b11110100101000:	sigmoid_prime = 18'b001010000001011000;
		14'b11110100101001:	sigmoid_prime = 18'b001010000010001001;
		14'b11110100101010:	sigmoid_prime = 18'b001010000010111010;
		14'b11110100101011:	sigmoid_prime = 18'b001010000011101011;
		14'b11110100101100:	sigmoid_prime = 18'b001010000100011100;
		14'b11110100101101:	sigmoid_prime = 18'b001010000101001110;
		14'b11110100101110:	sigmoid_prime = 18'b001010000101111111;
		14'b11110100101111:	sigmoid_prime = 18'b001010000110110000;
		14'b11110100110000:	sigmoid_prime = 18'b001010000111100001;
		14'b11110100110001:	sigmoid_prime = 18'b001010001000010010;
		14'b11110100110010:	sigmoid_prime = 18'b001010001001000011;
		14'b11110100110011:	sigmoid_prime = 18'b001010001001110100;
		14'b11110100110100:	sigmoid_prime = 18'b001010001010100101;
		14'b11110100110101:	sigmoid_prime = 18'b001010001011010110;
		14'b11110100110110:	sigmoid_prime = 18'b001010001100000111;
		14'b11110100110111:	sigmoid_prime = 18'b001010001100111000;
		14'b11110100111000:	sigmoid_prime = 18'b001010001101101010;
		14'b11110100111001:	sigmoid_prime = 18'b001010001110011011;
		14'b11110100111010:	sigmoid_prime = 18'b001010001111001100;
		14'b11110100111011:	sigmoid_prime = 18'b001010001111111101;
		14'b11110100111100:	sigmoid_prime = 18'b001010010000101110;
		14'b11110100111101:	sigmoid_prime = 18'b001010010001011111;
		14'b11110100111110:	sigmoid_prime = 18'b001010010010010001;
		14'b11110100111111:	sigmoid_prime = 18'b001010010011000010;
		14'b11110101000000:	sigmoid_prime = 18'b001010010011110011;
		14'b11110101000001:	sigmoid_prime = 18'b001010010100100100;
		14'b11110101000010:	sigmoid_prime = 18'b001010010101010101;
		14'b11110101000011:	sigmoid_prime = 18'b001010010110000110;
		14'b11110101000100:	sigmoid_prime = 18'b001010010110111000;
		14'b11110101000101:	sigmoid_prime = 18'b001010010111101001;
		14'b11110101000110:	sigmoid_prime = 18'b001010011000011010;
		14'b11110101000111:	sigmoid_prime = 18'b001010011001001011;
		14'b11110101001000:	sigmoid_prime = 18'b001010011001111101;
		14'b11110101001001:	sigmoid_prime = 18'b001010011010101110;
		14'b11110101001010:	sigmoid_prime = 18'b001010011011011111;
		14'b11110101001011:	sigmoid_prime = 18'b001010011100010000;
		14'b11110101001100:	sigmoid_prime = 18'b001010011101000001;
		14'b11110101001101:	sigmoid_prime = 18'b001010011101110011;
		14'b11110101001110:	sigmoid_prime = 18'b001010011110100100;
		14'b11110101001111:	sigmoid_prime = 18'b001010011111010101;
		14'b11110101010000:	sigmoid_prime = 18'b001010100000000110;
		14'b11110101010001:	sigmoid_prime = 18'b001010100000111000;
		14'b11110101010010:	sigmoid_prime = 18'b001010100001101001;
		14'b11110101010011:	sigmoid_prime = 18'b001010100010011010;
		14'b11110101010100:	sigmoid_prime = 18'b001010100011001011;
		14'b11110101010101:	sigmoid_prime = 18'b001010100011111101;
		14'b11110101010110:	sigmoid_prime = 18'b001010100100101110;
		14'b11110101010111:	sigmoid_prime = 18'b001010100101011111;
		14'b11110101011000:	sigmoid_prime = 18'b001010100110010000;
		14'b11110101011001:	sigmoid_prime = 18'b001010100111000010;
		14'b11110101011010:	sigmoid_prime = 18'b001010100111110011;
		14'b11110101011011:	sigmoid_prime = 18'b001010101000100100;
		14'b11110101011100:	sigmoid_prime = 18'b001010101001010110;
		14'b11110101011101:	sigmoid_prime = 18'b001010101010000111;
		14'b11110101011110:	sigmoid_prime = 18'b001010101010111000;
		14'b11110101011111:	sigmoid_prime = 18'b001010101011101001;
		14'b11110101100000:	sigmoid_prime = 18'b001010101100011011;
		14'b11110101100001:	sigmoid_prime = 18'b001010101101001100;
		14'b11110101100010:	sigmoid_prime = 18'b001010101101111101;
		14'b11110101100011:	sigmoid_prime = 18'b001010101110101110;
		14'b11110101100100:	sigmoid_prime = 18'b001010101111100000;
		14'b11110101100101:	sigmoid_prime = 18'b001010110000010001;
		14'b11110101100110:	sigmoid_prime = 18'b001010110001000010;
		14'b11110101100111:	sigmoid_prime = 18'b001010110001110011;
		14'b11110101101000:	sigmoid_prime = 18'b001010110010100101;
		14'b11110101101001:	sigmoid_prime = 18'b001010110011010110;
		14'b11110101101010:	sigmoid_prime = 18'b001010110100000111;
		14'b11110101101011:	sigmoid_prime = 18'b001010110100111000;
		14'b11110101101100:	sigmoid_prime = 18'b001010110101101010;
		14'b11110101101101:	sigmoid_prime = 18'b001010110110011011;
		14'b11110101101110:	sigmoid_prime = 18'b001010110111001100;
		14'b11110101101111:	sigmoid_prime = 18'b001010110111111101;
		14'b11110101110000:	sigmoid_prime = 18'b001010111000101111;
		14'b11110101110001:	sigmoid_prime = 18'b001010111001100000;
		14'b11110101110010:	sigmoid_prime = 18'b001010111010010001;
		14'b11110101110011:	sigmoid_prime = 18'b001010111011000010;
		14'b11110101110100:	sigmoid_prime = 18'b001010111011110100;
		14'b11110101110101:	sigmoid_prime = 18'b001010111100100101;
		14'b11110101110110:	sigmoid_prime = 18'b001010111101010110;
		14'b11110101110111:	sigmoid_prime = 18'b001010111110000111;
		14'b11110101111000:	sigmoid_prime = 18'b001010111110111000;
		14'b11110101111001:	sigmoid_prime = 18'b001010111111101010;
		14'b11110101111010:	sigmoid_prime = 18'b001011000000011011;
		14'b11110101111011:	sigmoid_prime = 18'b001011000001001100;
		14'b11110101111100:	sigmoid_prime = 18'b001011000001111101;
		14'b11110101111101:	sigmoid_prime = 18'b001011000010101110;
		14'b11110101111110:	sigmoid_prime = 18'b001011000011100000;
		14'b11110101111111:	sigmoid_prime = 18'b001011000100010001;
		14'b11110110000000:	sigmoid_prime = 18'b001011000101000010;
		14'b11110110000001:	sigmoid_prime = 18'b001011000101110011;
		14'b11110110000010:	sigmoid_prime = 18'b001011000110100100;
		14'b11110110000011:	sigmoid_prime = 18'b001011000111010101;
		14'b11110110000100:	sigmoid_prime = 18'b001011001000000110;
		14'b11110110000101:	sigmoid_prime = 18'b001011001000111000;
		14'b11110110000110:	sigmoid_prime = 18'b001011001001101001;
		14'b11110110000111:	sigmoid_prime = 18'b001011001010011010;
		14'b11110110001000:	sigmoid_prime = 18'b001011001011001011;
		14'b11110110001001:	sigmoid_prime = 18'b001011001011111100;
		14'b11110110001010:	sigmoid_prime = 18'b001011001100101101;
		14'b11110110001011:	sigmoid_prime = 18'b001011001101011110;
		14'b11110110001100:	sigmoid_prime = 18'b001011001110001111;
		14'b11110110001101:	sigmoid_prime = 18'b001011001111000000;
		14'b11110110001110:	sigmoid_prime = 18'b001011001111110001;
		14'b11110110001111:	sigmoid_prime = 18'b001011010000100010;
		14'b11110110010000:	sigmoid_prime = 18'b001011010001010011;
		14'b11110110010001:	sigmoid_prime = 18'b001011010010000100;
		14'b11110110010010:	sigmoid_prime = 18'b001011010010110101;
		14'b11110110010011:	sigmoid_prime = 18'b001011010011100110;
		14'b11110110010100:	sigmoid_prime = 18'b001011010100010111;
		14'b11110110010101:	sigmoid_prime = 18'b001011010101001000;
		14'b11110110010110:	sigmoid_prime = 18'b001011010101111001;
		14'b11110110010111:	sigmoid_prime = 18'b001011010110101010;
		14'b11110110011000:	sigmoid_prime = 18'b001011010111011011;
		14'b11110110011001:	sigmoid_prime = 18'b001011011000001100;
		14'b11110110011010:	sigmoid_prime = 18'b001011011000111101;
		14'b11110110011011:	sigmoid_prime = 18'b001011011001101110;
		14'b11110110011100:	sigmoid_prime = 18'b001011011010011111;
		14'b11110110011101:	sigmoid_prime = 18'b001011011011010000;
		14'b11110110011110:	sigmoid_prime = 18'b001011011100000001;
		14'b11110110011111:	sigmoid_prime = 18'b001011011100110001;
		14'b11110110100000:	sigmoid_prime = 18'b001011011101100010;
		14'b11110110100001:	sigmoid_prime = 18'b001011011110010011;
		14'b11110110100010:	sigmoid_prime = 18'b001011011111000100;
		14'b11110110100011:	sigmoid_prime = 18'b001011011111110101;
		14'b11110110100100:	sigmoid_prime = 18'b001011100000100101;
		14'b11110110100101:	sigmoid_prime = 18'b001011100001010110;
		14'b11110110100110:	sigmoid_prime = 18'b001011100010000111;
		14'b11110110100111:	sigmoid_prime = 18'b001011100010111000;
		14'b11110110101000:	sigmoid_prime = 18'b001011100011101000;
		14'b11110110101001:	sigmoid_prime = 18'b001011100100011001;
		14'b11110110101010:	sigmoid_prime = 18'b001011100101001010;
		14'b11110110101011:	sigmoid_prime = 18'b001011100101111011;
		14'b11110110101100:	sigmoid_prime = 18'b001011100110101011;
		14'b11110110101101:	sigmoid_prime = 18'b001011100111011100;
		14'b11110110101110:	sigmoid_prime = 18'b001011101000001101;
		14'b11110110101111:	sigmoid_prime = 18'b001011101000111101;
		14'b11110110110000:	sigmoid_prime = 18'b001011101001101110;
		14'b11110110110001:	sigmoid_prime = 18'b001011101010011110;
		14'b11110110110010:	sigmoid_prime = 18'b001011101011001111;
		14'b11110110110011:	sigmoid_prime = 18'b001011101011111111;
		14'b11110110110100:	sigmoid_prime = 18'b001011101100110000;
		14'b11110110110101:	sigmoid_prime = 18'b001011101101100001;
		14'b11110110110110:	sigmoid_prime = 18'b001011101110010001;
		14'b11110110110111:	sigmoid_prime = 18'b001011101111000001;
		14'b11110110111000:	sigmoid_prime = 18'b001011101111110010;
		14'b11110110111001:	sigmoid_prime = 18'b001011110000100010;
		14'b11110110111010:	sigmoid_prime = 18'b001011110001010011;
		14'b11110110111011:	sigmoid_prime = 18'b001011110010000011;
		14'b11110110111100:	sigmoid_prime = 18'b001011110010110100;
		14'b11110110111101:	sigmoid_prime = 18'b001011110011100100;
		14'b11110110111110:	sigmoid_prime = 18'b001011110100010100;
		14'b11110110111111:	sigmoid_prime = 18'b001011110101000101;
		14'b11110111000000:	sigmoid_prime = 18'b001011110101110101;
		14'b11110111000001:	sigmoid_prime = 18'b001011110110100101;
		14'b11110111000010:	sigmoid_prime = 18'b001011110111010110;
		14'b11110111000011:	sigmoid_prime = 18'b001011111000000110;
		14'b11110111000100:	sigmoid_prime = 18'b001011111000110110;
		14'b11110111000101:	sigmoid_prime = 18'b001011111001100110;
		14'b11110111000110:	sigmoid_prime = 18'b001011111010010110;
		14'b11110111000111:	sigmoid_prime = 18'b001011111011000111;
		14'b11110111001000:	sigmoid_prime = 18'b001011111011110111;
		14'b11110111001001:	sigmoid_prime = 18'b001011111100100111;
		14'b11110111001010:	sigmoid_prime = 18'b001011111101010111;
		14'b11110111001011:	sigmoid_prime = 18'b001011111110000111;
		14'b11110111001100:	sigmoid_prime = 18'b001011111110110111;
		14'b11110111001101:	sigmoid_prime = 18'b001011111111100111;
		14'b11110111001110:	sigmoid_prime = 18'b001100000000010111;
		14'b11110111001111:	sigmoid_prime = 18'b001100000001000111;
		14'b11110111010000:	sigmoid_prime = 18'b001100000001110111;
		14'b11110111010001:	sigmoid_prime = 18'b001100000010100111;
		14'b11110111010010:	sigmoid_prime = 18'b001100000011010111;
		14'b11110111010011:	sigmoid_prime = 18'b001100000100000111;
		14'b11110111010100:	sigmoid_prime = 18'b001100000100110110;
		14'b11110111010101:	sigmoid_prime = 18'b001100000101100110;
		14'b11110111010110:	sigmoid_prime = 18'b001100000110010110;
		14'b11110111010111:	sigmoid_prime = 18'b001100000111000110;
		14'b11110111011000:	sigmoid_prime = 18'b001100000111110110;
		14'b11110111011001:	sigmoid_prime = 18'b001100001000100101;
		14'b11110111011010:	sigmoid_prime = 18'b001100001001010101;
		14'b11110111011011:	sigmoid_prime = 18'b001100001010000101;
		14'b11110111011100:	sigmoid_prime = 18'b001100001010110100;
		14'b11110111011101:	sigmoid_prime = 18'b001100001011100100;
		14'b11110111011110:	sigmoid_prime = 18'b001100001100010100;
		14'b11110111011111:	sigmoid_prime = 18'b001100001101000011;
		14'b11110111100000:	sigmoid_prime = 18'b001100001101110011;
		14'b11110111100001:	sigmoid_prime = 18'b001100001110100010;
		14'b11110111100010:	sigmoid_prime = 18'b001100001111010010;
		14'b11110111100011:	sigmoid_prime = 18'b001100010000000001;
		14'b11110111100100:	sigmoid_prime = 18'b001100010000110001;
		14'b11110111100101:	sigmoid_prime = 18'b001100010001100000;
		14'b11110111100110:	sigmoid_prime = 18'b001100010010001111;
		14'b11110111100111:	sigmoid_prime = 18'b001100010010111111;
		14'b11110111101000:	sigmoid_prime = 18'b001100010011101110;
		14'b11110111101001:	sigmoid_prime = 18'b001100010100011101;
		14'b11110111101010:	sigmoid_prime = 18'b001100010101001101;
		14'b11110111101011:	sigmoid_prime = 18'b001100010101111100;
		14'b11110111101100:	sigmoid_prime = 18'b001100010110101011;
		14'b11110111101101:	sigmoid_prime = 18'b001100010111011010;
		14'b11110111101110:	sigmoid_prime = 18'b001100011000001001;
		14'b11110111101111:	sigmoid_prime = 18'b001100011000111000;
		14'b11110111110000:	sigmoid_prime = 18'b001100011001100111;
		14'b11110111110001:	sigmoid_prime = 18'b001100011010010111;
		14'b11110111110010:	sigmoid_prime = 18'b001100011011000110;
		14'b11110111110011:	sigmoid_prime = 18'b001100011011110100;
		14'b11110111110100:	sigmoid_prime = 18'b001100011100100011;
		14'b11110111110101:	sigmoid_prime = 18'b001100011101010010;
		14'b11110111110110:	sigmoid_prime = 18'b001100011110000001;
		14'b11110111110111:	sigmoid_prime = 18'b001100011110110000;
		14'b11110111111000:	sigmoid_prime = 18'b001100011111011111;
		14'b11110111111001:	sigmoid_prime = 18'b001100100000001110;
		14'b11110111111010:	sigmoid_prime = 18'b001100100000111100;
		14'b11110111111011:	sigmoid_prime = 18'b001100100001101011;
		14'b11110111111100:	sigmoid_prime = 18'b001100100010011010;
		14'b11110111111101:	sigmoid_prime = 18'b001100100011001000;
		14'b11110111111110:	sigmoid_prime = 18'b001100100011110111;
		14'b11110111111111:	sigmoid_prime = 18'b001100100100100110;
		14'b11111000000000:	sigmoid_prime = 18'b001100100101010100;
		14'b11111000000001:	sigmoid_prime = 18'b001100100110000011;
		14'b11111000000010:	sigmoid_prime = 18'b001100100110110001;
		14'b11111000000011:	sigmoid_prime = 18'b001100100111100000;
		14'b11111000000100:	sigmoid_prime = 18'b001100101000001110;
		14'b11111000000101:	sigmoid_prime = 18'b001100101000111100;
		14'b11111000000110:	sigmoid_prime = 18'b001100101001101011;
		14'b11111000000111:	sigmoid_prime = 18'b001100101010011001;
		14'b11111000001000:	sigmoid_prime = 18'b001100101011000111;
		14'b11111000001001:	sigmoid_prime = 18'b001100101011110101;
		14'b11111000001010:	sigmoid_prime = 18'b001100101100100100;
		14'b11111000001011:	sigmoid_prime = 18'b001100101101010010;
		14'b11111000001100:	sigmoid_prime = 18'b001100101110000000;
		14'b11111000001101:	sigmoid_prime = 18'b001100101110101110;
		14'b11111000001110:	sigmoid_prime = 18'b001100101111011100;
		14'b11111000001111:	sigmoid_prime = 18'b001100110000001010;
		14'b11111000010000:	sigmoid_prime = 18'b001100110000111000;
		14'b11111000010001:	sigmoid_prime = 18'b001100110001100110;
		14'b11111000010010:	sigmoid_prime = 18'b001100110010010100;
		14'b11111000010011:	sigmoid_prime = 18'b001100110011000001;
		14'b11111000010100:	sigmoid_prime = 18'b001100110011101111;
		14'b11111000010101:	sigmoid_prime = 18'b001100110100011101;
		14'b11111000010110:	sigmoid_prime = 18'b001100110101001011;
		14'b11111000010111:	sigmoid_prime = 18'b001100110101111000;
		14'b11111000011000:	sigmoid_prime = 18'b001100110110100110;
		14'b11111000011001:	sigmoid_prime = 18'b001100110111010011;
		14'b11111000011010:	sigmoid_prime = 18'b001100111000000001;
		14'b11111000011011:	sigmoid_prime = 18'b001100111000101110;
		14'b11111000011100:	sigmoid_prime = 18'b001100111001011100;
		14'b11111000011101:	sigmoid_prime = 18'b001100111010001001;
		14'b11111000011110:	sigmoid_prime = 18'b001100111010110111;
		14'b11111000011111:	sigmoid_prime = 18'b001100111011100100;
		14'b11111000100000:	sigmoid_prime = 18'b001100111100010001;
		14'b11111000100001:	sigmoid_prime = 18'b001100111100111111;
		14'b11111000100010:	sigmoid_prime = 18'b001100111101101100;
		14'b11111000100011:	sigmoid_prime = 18'b001100111110011001;
		14'b11111000100100:	sigmoid_prime = 18'b001100111111000110;
		14'b11111000100101:	sigmoid_prime = 18'b001100111111110011;
		14'b11111000100110:	sigmoid_prime = 18'b001101000000100000;
		14'b11111000100111:	sigmoid_prime = 18'b001101000001001101;
		14'b11111000101000:	sigmoid_prime = 18'b001101000001111010;
		14'b11111000101001:	sigmoid_prime = 18'b001101000010100111;
		14'b11111000101010:	sigmoid_prime = 18'b001101000011010100;
		14'b11111000101011:	sigmoid_prime = 18'b001101000100000001;
		14'b11111000101100:	sigmoid_prime = 18'b001101000100101101;
		14'b11111000101101:	sigmoid_prime = 18'b001101000101011010;
		14'b11111000101110:	sigmoid_prime = 18'b001101000110000111;
		14'b11111000101111:	sigmoid_prime = 18'b001101000110110011;
		14'b11111000110000:	sigmoid_prime = 18'b001101000111100000;
		14'b11111000110001:	sigmoid_prime = 18'b001101001000001100;
		14'b11111000110010:	sigmoid_prime = 18'b001101001000111001;
		14'b11111000110011:	sigmoid_prime = 18'b001101001001100101;
		14'b11111000110100:	sigmoid_prime = 18'b001101001010010010;
		14'b11111000110101:	sigmoid_prime = 18'b001101001010111110;
		14'b11111000110110:	sigmoid_prime = 18'b001101001011101010;
		14'b11111000110111:	sigmoid_prime = 18'b001101001100010111;
		14'b11111000111000:	sigmoid_prime = 18'b001101001101000011;
		14'b11111000111001:	sigmoid_prime = 18'b001101001101101111;
		14'b11111000111010:	sigmoid_prime = 18'b001101001110011011;
		14'b11111000111011:	sigmoid_prime = 18'b001101001111000111;
		14'b11111000111100:	sigmoid_prime = 18'b001101001111110011;
		14'b11111000111101:	sigmoid_prime = 18'b001101010000011111;
		14'b11111000111110:	sigmoid_prime = 18'b001101010001001011;
		14'b11111000111111:	sigmoid_prime = 18'b001101010001110111;
		14'b11111001000000:	sigmoid_prime = 18'b001101010010100010;
		14'b11111001000001:	sigmoid_prime = 18'b001101010011001110;
		14'b11111001000010:	sigmoid_prime = 18'b001101010011111010;
		14'b11111001000011:	sigmoid_prime = 18'b001101010100100101;
		14'b11111001000100:	sigmoid_prime = 18'b001101010101010001;
		14'b11111001000101:	sigmoid_prime = 18'b001101010101111101;
		14'b11111001000110:	sigmoid_prime = 18'b001101010110101000;
		14'b11111001000111:	sigmoid_prime = 18'b001101010111010011;
		14'b11111001001000:	sigmoid_prime = 18'b001101010111111111;
		14'b11111001001001:	sigmoid_prime = 18'b001101011000101010;
		14'b11111001001010:	sigmoid_prime = 18'b001101011001010101;
		14'b11111001001011:	sigmoid_prime = 18'b001101011010000001;
		14'b11111001001100:	sigmoid_prime = 18'b001101011010101100;
		14'b11111001001101:	sigmoid_prime = 18'b001101011011010111;
		14'b11111001001110:	sigmoid_prime = 18'b001101011100000010;
		14'b11111001001111:	sigmoid_prime = 18'b001101011100101101;
		14'b11111001010000:	sigmoid_prime = 18'b001101011101011000;
		14'b11111001010001:	sigmoid_prime = 18'b001101011110000011;
		14'b11111001010010:	sigmoid_prime = 18'b001101011110101101;
		14'b11111001010011:	sigmoid_prime = 18'b001101011111011000;
		14'b11111001010100:	sigmoid_prime = 18'b001101100000000011;
		14'b11111001010101:	sigmoid_prime = 18'b001101100000101110;
		14'b11111001010110:	sigmoid_prime = 18'b001101100001011000;
		14'b11111001010111:	sigmoid_prime = 18'b001101100010000011;
		14'b11111001011000:	sigmoid_prime = 18'b001101100010101101;
		14'b11111001011001:	sigmoid_prime = 18'b001101100011011000;
		14'b11111001011010:	sigmoid_prime = 18'b001101100100000010;
		14'b11111001011011:	sigmoid_prime = 18'b001101100100101100;
		14'b11111001011100:	sigmoid_prime = 18'b001101100101010111;
		14'b11111001011101:	sigmoid_prime = 18'b001101100110000001;
		14'b11111001011110:	sigmoid_prime = 18'b001101100110101011;
		14'b11111001011111:	sigmoid_prime = 18'b001101100111010101;
		14'b11111001100000:	sigmoid_prime = 18'b001101100111111111;
		14'b11111001100001:	sigmoid_prime = 18'b001101101000101001;
		14'b11111001100010:	sigmoid_prime = 18'b001101101001010011;
		14'b11111001100011:	sigmoid_prime = 18'b001101101001111101;
		14'b11111001100100:	sigmoid_prime = 18'b001101101010100111;
		14'b11111001100101:	sigmoid_prime = 18'b001101101011010000;
		14'b11111001100110:	sigmoid_prime = 18'b001101101011111010;
		14'b11111001100111:	sigmoid_prime = 18'b001101101100100100;
		14'b11111001101000:	sigmoid_prime = 18'b001101101101001101;
		14'b11111001101001:	sigmoid_prime = 18'b001101101101110111;
		14'b11111001101010:	sigmoid_prime = 18'b001101101110100000;
		14'b11111001101011:	sigmoid_prime = 18'b001101101111001001;
		14'b11111001101100:	sigmoid_prime = 18'b001101101111110011;
		14'b11111001101101:	sigmoid_prime = 18'b001101110000011100;
		14'b11111001101110:	sigmoid_prime = 18'b001101110001000101;
		14'b11111001101111:	sigmoid_prime = 18'b001101110001101110;
		14'b11111001110000:	sigmoid_prime = 18'b001101110010010111;
		14'b11111001110001:	sigmoid_prime = 18'b001101110011000000;
		14'b11111001110010:	sigmoid_prime = 18'b001101110011101001;
		14'b11111001110011:	sigmoid_prime = 18'b001101110100010010;
		14'b11111001110100:	sigmoid_prime = 18'b001101110100111011;
		14'b11111001110101:	sigmoid_prime = 18'b001101110101100100;
		14'b11111001110110:	sigmoid_prime = 18'b001101110110001100;
		14'b11111001110111:	sigmoid_prime = 18'b001101110110110101;
		14'b11111001111000:	sigmoid_prime = 18'b001101110111011101;
		14'b11111001111001:	sigmoid_prime = 18'b001101111000000110;
		14'b11111001111010:	sigmoid_prime = 18'b001101111000101110;
		14'b11111001111011:	sigmoid_prime = 18'b001101111001010111;
		14'b11111001111100:	sigmoid_prime = 18'b001101111001111111;
		14'b11111001111101:	sigmoid_prime = 18'b001101111010100111;
		14'b11111001111110:	sigmoid_prime = 18'b001101111011001111;
		14'b11111001111111:	sigmoid_prime = 18'b001101111011110111;
		14'b11111010000000:	sigmoid_prime = 18'b001101111100011111;
		14'b11111010000001:	sigmoid_prime = 18'b001101111101000111;
		14'b11111010000010:	sigmoid_prime = 18'b001101111101101111;
		14'b11111010000011:	sigmoid_prime = 18'b001101111110010111;
		14'b11111010000100:	sigmoid_prime = 18'b001101111110111111;
		14'b11111010000101:	sigmoid_prime = 18'b001101111111100110;
		14'b11111010000110:	sigmoid_prime = 18'b001110000000001110;
		14'b11111010000111:	sigmoid_prime = 18'b001110000000110110;
		14'b11111010001000:	sigmoid_prime = 18'b001110000001011101;
		14'b11111010001001:	sigmoid_prime = 18'b001110000010000100;
		14'b11111010001010:	sigmoid_prime = 18'b001110000010101100;
		14'b11111010001011:	sigmoid_prime = 18'b001110000011010011;
		14'b11111010001100:	sigmoid_prime = 18'b001110000011111010;
		14'b11111010001101:	sigmoid_prime = 18'b001110000100100001;
		14'b11111010001110:	sigmoid_prime = 18'b001110000101001000;
		14'b11111010001111:	sigmoid_prime = 18'b001110000101101111;
		14'b11111010010000:	sigmoid_prime = 18'b001110000110010110;
		14'b11111010010001:	sigmoid_prime = 18'b001110000110111101;
		14'b11111010010010:	sigmoid_prime = 18'b001110000111100100;
		14'b11111010010011:	sigmoid_prime = 18'b001110001000001011;
		14'b11111010010100:	sigmoid_prime = 18'b001110001000110001;
		14'b11111010010101:	sigmoid_prime = 18'b001110001001011000;
		14'b11111010010110:	sigmoid_prime = 18'b001110001001111110;
		14'b11111010010111:	sigmoid_prime = 18'b001110001010100101;
		14'b11111010011000:	sigmoid_prime = 18'b001110001011001011;
		14'b11111010011001:	sigmoid_prime = 18'b001110001011110001;
		14'b11111010011010:	sigmoid_prime = 18'b001110001100010111;
		14'b11111010011011:	sigmoid_prime = 18'b001110001100111110;
		14'b11111010011100:	sigmoid_prime = 18'b001110001101100100;
		14'b11111010011101:	sigmoid_prime = 18'b001110001110001010;
		14'b11111010011110:	sigmoid_prime = 18'b001110001110101111;
		14'b11111010011111:	sigmoid_prime = 18'b001110001111010101;
		14'b11111010100000:	sigmoid_prime = 18'b001110001111111011;
		14'b11111010100001:	sigmoid_prime = 18'b001110010000100001;
		14'b11111010100010:	sigmoid_prime = 18'b001110010001000110;
		14'b11111010100011:	sigmoid_prime = 18'b001110010001101100;
		14'b11111010100100:	sigmoid_prime = 18'b001110010010010001;
		14'b11111010100101:	sigmoid_prime = 18'b001110010010110111;
		14'b11111010100110:	sigmoid_prime = 18'b001110010011011100;
		14'b11111010100111:	sigmoid_prime = 18'b001110010100000001;
		14'b11111010101000:	sigmoid_prime = 18'b001110010100100110;
		14'b11111010101001:	sigmoid_prime = 18'b001110010101001011;
		14'b11111010101010:	sigmoid_prime = 18'b001110010101110000;
		14'b11111010101011:	sigmoid_prime = 18'b001110010110010101;
		14'b11111010101100:	sigmoid_prime = 18'b001110010110111010;
		14'b11111010101101:	sigmoid_prime = 18'b001110010111011111;
		14'b11111010101110:	sigmoid_prime = 18'b001110011000000100;
		14'b11111010101111:	sigmoid_prime = 18'b001110011000101000;
		14'b11111010110000:	sigmoid_prime = 18'b001110011001001101;
		14'b11111010110001:	sigmoid_prime = 18'b001110011001110001;
		14'b11111010110010:	sigmoid_prime = 18'b001110011010010110;
		14'b11111010110011:	sigmoid_prime = 18'b001110011010111010;
		14'b11111010110100:	sigmoid_prime = 18'b001110011011011110;
		14'b11111010110101:	sigmoid_prime = 18'b001110011100000010;
		14'b11111010110110:	sigmoid_prime = 18'b001110011100100110;
		14'b11111010110111:	sigmoid_prime = 18'b001110011101001010;
		14'b11111010111000:	sigmoid_prime = 18'b001110011101101110;
		14'b11111010111001:	sigmoid_prime = 18'b001110011110010010;
		14'b11111010111010:	sigmoid_prime = 18'b001110011110110110;
		14'b11111010111011:	sigmoid_prime = 18'b001110011111011001;
		14'b11111010111100:	sigmoid_prime = 18'b001110011111111101;
		14'b11111010111101:	sigmoid_prime = 18'b001110100000100000;
		14'b11111010111110:	sigmoid_prime = 18'b001110100001000100;
		14'b11111010111111:	sigmoid_prime = 18'b001110100001100111;
		14'b11111011000000:	sigmoid_prime = 18'b001110100010001010;
		14'b11111011000001:	sigmoid_prime = 18'b001110100010101101;
		14'b11111011000010:	sigmoid_prime = 18'b001110100011010000;
		14'b11111011000011:	sigmoid_prime = 18'b001110100011110011;
		14'b11111011000100:	sigmoid_prime = 18'b001110100100010110;
		14'b11111011000101:	sigmoid_prime = 18'b001110100100111001;
		14'b11111011000110:	sigmoid_prime = 18'b001110100101011100;
		14'b11111011000111:	sigmoid_prime = 18'b001110100101111111;
		14'b11111011001000:	sigmoid_prime = 18'b001110100110100001;
		14'b11111011001001:	sigmoid_prime = 18'b001110100111000100;
		14'b11111011001010:	sigmoid_prime = 18'b001110100111100110;
		14'b11111011001011:	sigmoid_prime = 18'b001110101000001000;
		14'b11111011001100:	sigmoid_prime = 18'b001110101000101011;
		14'b11111011001101:	sigmoid_prime = 18'b001110101001001101;
		14'b11111011001110:	sigmoid_prime = 18'b001110101001101111;
		14'b11111011001111:	sigmoid_prime = 18'b001110101010010001;
		14'b11111011010000:	sigmoid_prime = 18'b001110101010110011;
		14'b11111011010001:	sigmoid_prime = 18'b001110101011010100;
		14'b11111011010010:	sigmoid_prime = 18'b001110101011110110;
		14'b11111011010011:	sigmoid_prime = 18'b001110101100011000;
		14'b11111011010100:	sigmoid_prime = 18'b001110101100111001;
		14'b11111011010101:	sigmoid_prime = 18'b001110101101011011;
		14'b11111011010110:	sigmoid_prime = 18'b001110101101111100;
		14'b11111011010111:	sigmoid_prime = 18'b001110101110011110;
		14'b11111011011000:	sigmoid_prime = 18'b001110101110111111;
		14'b11111011011001:	sigmoid_prime = 18'b001110101111100000;
		14'b11111011011010:	sigmoid_prime = 18'b001110110000000001;
		14'b11111011011011:	sigmoid_prime = 18'b001110110000100010;
		14'b11111011011100:	sigmoid_prime = 18'b001110110001000011;
		14'b11111011011101:	sigmoid_prime = 18'b001110110001100011;
		14'b11111011011110:	sigmoid_prime = 18'b001110110010000100;
		14'b11111011011111:	sigmoid_prime = 18'b001110110010100101;
		14'b11111011100000:	sigmoid_prime = 18'b001110110011000101;
		14'b11111011100001:	sigmoid_prime = 18'b001110110011100110;
		14'b11111011100010:	sigmoid_prime = 18'b001110110100000110;
		14'b11111011100011:	sigmoid_prime = 18'b001110110100100110;
		14'b11111011100100:	sigmoid_prime = 18'b001110110101000110;
		14'b11111011100101:	sigmoid_prime = 18'b001110110101100110;
		14'b11111011100110:	sigmoid_prime = 18'b001110110110000110;
		14'b11111011100111:	sigmoid_prime = 18'b001110110110100110;
		14'b11111011101000:	sigmoid_prime = 18'b001110110111000110;
		14'b11111011101001:	sigmoid_prime = 18'b001110110111100101;
		14'b11111011101010:	sigmoid_prime = 18'b001110111000000101;
		14'b11111011101011:	sigmoid_prime = 18'b001110111000100101;
		14'b11111011101100:	sigmoid_prime = 18'b001110111001000100;
		14'b11111011101101:	sigmoid_prime = 18'b001110111001100011;
		14'b11111011101110:	sigmoid_prime = 18'b001110111010000010;
		14'b11111011101111:	sigmoid_prime = 18'b001110111010100010;
		14'b11111011110000:	sigmoid_prime = 18'b001110111011000001;
		14'b11111011110001:	sigmoid_prime = 18'b001110111011100000;
		14'b11111011110010:	sigmoid_prime = 18'b001110111011111110;
		14'b11111011110011:	sigmoid_prime = 18'b001110111100011101;
		14'b11111011110100:	sigmoid_prime = 18'b001110111100111100;
		14'b11111011110101:	sigmoid_prime = 18'b001110111101011010;
		14'b11111011110110:	sigmoid_prime = 18'b001110111101111001;
		14'b11111011110111:	sigmoid_prime = 18'b001110111110010111;
		14'b11111011111000:	sigmoid_prime = 18'b001110111110110101;
		14'b11111011111001:	sigmoid_prime = 18'b001110111111010100;
		14'b11111011111010:	sigmoid_prime = 18'b001110111111110010;
		14'b11111011111011:	sigmoid_prime = 18'b001111000000010000;
		14'b11111011111100:	sigmoid_prime = 18'b001111000000101110;
		14'b11111011111101:	sigmoid_prime = 18'b001111000001001011;
		14'b11111011111110:	sigmoid_prime = 18'b001111000001101001;
		14'b11111011111111:	sigmoid_prime = 18'b001111000010000111;
		14'b11111100000000:	sigmoid_prime = 18'b001111000010100100;
		14'b11111100000001:	sigmoid_prime = 18'b001111000011000010;
		14'b11111100000010:	sigmoid_prime = 18'b001111000011011111;
		14'b11111100000011:	sigmoid_prime = 18'b001111000011111100;
		14'b11111100000100:	sigmoid_prime = 18'b001111000100011001;
		14'b11111100000101:	sigmoid_prime = 18'b001111000100110110;
		14'b11111100000110:	sigmoid_prime = 18'b001111000101010011;
		14'b11111100000111:	sigmoid_prime = 18'b001111000101110000;
		14'b11111100001000:	sigmoid_prime = 18'b001111000110001101;
		14'b11111100001001:	sigmoid_prime = 18'b001111000110101010;
		14'b11111100001010:	sigmoid_prime = 18'b001111000111000110;
		14'b11111100001011:	sigmoid_prime = 18'b001111000111100011;
		14'b11111100001100:	sigmoid_prime = 18'b001111000111111111;
		14'b11111100001101:	sigmoid_prime = 18'b001111001000011011;
		14'b11111100001110:	sigmoid_prime = 18'b001111001000110111;
		14'b11111100001111:	sigmoid_prime = 18'b001111001001010011;
		14'b11111100010000:	sigmoid_prime = 18'b001111001001101111;
		14'b11111100010001:	sigmoid_prime = 18'b001111001010001011;
		14'b11111100010010:	sigmoid_prime = 18'b001111001010100111;
		14'b11111100010011:	sigmoid_prime = 18'b001111001011000011;
		14'b11111100010100:	sigmoid_prime = 18'b001111001011011110;
		14'b11111100010101:	sigmoid_prime = 18'b001111001011111010;
		14'b11111100010110:	sigmoid_prime = 18'b001111001100010101;
		14'b11111100010111:	sigmoid_prime = 18'b001111001100110000;
		14'b11111100011000:	sigmoid_prime = 18'b001111001101001011;
		14'b11111100011001:	sigmoid_prime = 18'b001111001101100110;
		14'b11111100011010:	sigmoid_prime = 18'b001111001110000001;
		14'b11111100011011:	sigmoid_prime = 18'b001111001110011100;
		14'b11111100011100:	sigmoid_prime = 18'b001111001110110111;
		14'b11111100011101:	sigmoid_prime = 18'b001111001111010010;
		14'b11111100011110:	sigmoid_prime = 18'b001111001111101100;
		14'b11111100011111:	sigmoid_prime = 18'b001111010000000111;
		14'b11111100100000:	sigmoid_prime = 18'b001111010000100001;
		14'b11111100100001:	sigmoid_prime = 18'b001111010000111011;
		14'b11111100100010:	sigmoid_prime = 18'b001111010001010101;
		14'b11111100100011:	sigmoid_prime = 18'b001111010001101111;
		14'b11111100100100:	sigmoid_prime = 18'b001111010010001001;
		14'b11111100100101:	sigmoid_prime = 18'b001111010010100011;
		14'b11111100100110:	sigmoid_prime = 18'b001111010010111101;
		14'b11111100100111:	sigmoid_prime = 18'b001111010011010110;
		14'b11111100101000:	sigmoid_prime = 18'b001111010011110000;
		14'b11111100101001:	sigmoid_prime = 18'b001111010100001001;
		14'b11111100101010:	sigmoid_prime = 18'b001111010100100011;
		14'b11111100101011:	sigmoid_prime = 18'b001111010100111100;
		14'b11111100101100:	sigmoid_prime = 18'b001111010101010101;
		14'b11111100101101:	sigmoid_prime = 18'b001111010101101110;
		14'b11111100101110:	sigmoid_prime = 18'b001111010110000111;
		14'b11111100101111:	sigmoid_prime = 18'b001111010110100000;
		14'b11111100110000:	sigmoid_prime = 18'b001111010110111000;
		14'b11111100110001:	sigmoid_prime = 18'b001111010111010001;
		14'b11111100110010:	sigmoid_prime = 18'b001111010111101001;
		14'b11111100110011:	sigmoid_prime = 18'b001111011000000010;
		14'b11111100110100:	sigmoid_prime = 18'b001111011000011010;
		14'b11111100110101:	sigmoid_prime = 18'b001111011000110010;
		14'b11111100110110:	sigmoid_prime = 18'b001111011001001010;
		14'b11111100110111:	sigmoid_prime = 18'b001111011001100010;
		14'b11111100111000:	sigmoid_prime = 18'b001111011001111010;
		14'b11111100111001:	sigmoid_prime = 18'b001111011010010001;
		14'b11111100111010:	sigmoid_prime = 18'b001111011010101001;
		14'b11111100111011:	sigmoid_prime = 18'b001111011011000001;
		14'b11111100111100:	sigmoid_prime = 18'b001111011011011000;
		14'b11111100111101:	sigmoid_prime = 18'b001111011011101111;
		14'b11111100111110:	sigmoid_prime = 18'b001111011100000110;
		14'b11111100111111:	sigmoid_prime = 18'b001111011100011101;
		14'b11111101000000:	sigmoid_prime = 18'b001111011100110100;
		14'b11111101000001:	sigmoid_prime = 18'b001111011101001011;
		14'b11111101000010:	sigmoid_prime = 18'b001111011101100010;
		14'b11111101000011:	sigmoid_prime = 18'b001111011101111001;
		14'b11111101000100:	sigmoid_prime = 18'b001111011110001111;
		14'b11111101000101:	sigmoid_prime = 18'b001111011110100110;
		14'b11111101000110:	sigmoid_prime = 18'b001111011110111100;
		14'b11111101000111:	sigmoid_prime = 18'b001111011111010010;
		14'b11111101001000:	sigmoid_prime = 18'b001111011111101000;
		14'b11111101001001:	sigmoid_prime = 18'b001111011111111110;
		14'b11111101001010:	sigmoid_prime = 18'b001111100000010100;
		14'b11111101001011:	sigmoid_prime = 18'b001111100000101010;
		14'b11111101001100:	sigmoid_prime = 18'b001111100000111111;
		14'b11111101001101:	sigmoid_prime = 18'b001111100001010101;
		14'b11111101001110:	sigmoid_prime = 18'b001111100001101010;
		14'b11111101001111:	sigmoid_prime = 18'b001111100010000000;
		14'b11111101010000:	sigmoid_prime = 18'b001111100010010101;
		14'b11111101010001:	sigmoid_prime = 18'b001111100010101010;
		14'b11111101010010:	sigmoid_prime = 18'b001111100010111111;
		14'b11111101010011:	sigmoid_prime = 18'b001111100011010100;
		14'b11111101010100:	sigmoid_prime = 18'b001111100011101001;
		14'b11111101010101:	sigmoid_prime = 18'b001111100011111101;
		14'b11111101010110:	sigmoid_prime = 18'b001111100100010010;
		14'b11111101010111:	sigmoid_prime = 18'b001111100100100110;
		14'b11111101011000:	sigmoid_prime = 18'b001111100100111011;
		14'b11111101011001:	sigmoid_prime = 18'b001111100101001111;
		14'b11111101011010:	sigmoid_prime = 18'b001111100101100011;
		14'b11111101011011:	sigmoid_prime = 18'b001111100101110111;
		14'b11111101011100:	sigmoid_prime = 18'b001111100110001011;
		14'b11111101011101:	sigmoid_prime = 18'b001111100110011111;
		14'b11111101011110:	sigmoid_prime = 18'b001111100110110010;
		14'b11111101011111:	sigmoid_prime = 18'b001111100111000110;
		14'b11111101100000:	sigmoid_prime = 18'b001111100111011001;
		14'b11111101100001:	sigmoid_prime = 18'b001111100111101100;
		14'b11111101100010:	sigmoid_prime = 18'b001111101000000000;
		14'b11111101100011:	sigmoid_prime = 18'b001111101000010011;
		14'b11111101100100:	sigmoid_prime = 18'b001111101000100110;
		14'b11111101100101:	sigmoid_prime = 18'b001111101000111001;
		14'b11111101100110:	sigmoid_prime = 18'b001111101001001011;
		14'b11111101100111:	sigmoid_prime = 18'b001111101001011110;
		14'b11111101101000:	sigmoid_prime = 18'b001111101001110000;
		14'b11111101101001:	sigmoid_prime = 18'b001111101010000011;
		14'b11111101101010:	sigmoid_prime = 18'b001111101010010101;
		14'b11111101101011:	sigmoid_prime = 18'b001111101010100111;
		14'b11111101101100:	sigmoid_prime = 18'b001111101010111001;
		14'b11111101101101:	sigmoid_prime = 18'b001111101011001011;
		14'b11111101101110:	sigmoid_prime = 18'b001111101011011101;
		14'b11111101101111:	sigmoid_prime = 18'b001111101011101111;
		14'b11111101110000:	sigmoid_prime = 18'b001111101100000000;
		14'b11111101110001:	sigmoid_prime = 18'b001111101100010010;
		14'b11111101110010:	sigmoid_prime = 18'b001111101100100011;
		14'b11111101110011:	sigmoid_prime = 18'b001111101100110100;
		14'b11111101110100:	sigmoid_prime = 18'b001111101101000110;
		14'b11111101110101:	sigmoid_prime = 18'b001111101101010111;
		14'b11111101110110:	sigmoid_prime = 18'b001111101101101000;
		14'b11111101110111:	sigmoid_prime = 18'b001111101101111000;
		14'b11111101111000:	sigmoid_prime = 18'b001111101110001001;
		14'b11111101111001:	sigmoid_prime = 18'b001111101110011010;
		14'b11111101111010:	sigmoid_prime = 18'b001111101110101010;
		14'b11111101111011:	sigmoid_prime = 18'b001111101110111010;
		14'b11111101111100:	sigmoid_prime = 18'b001111101111001010;
		14'b11111101111101:	sigmoid_prime = 18'b001111101111011011;
		14'b11111101111110:	sigmoid_prime = 18'b001111101111101010;
		14'b11111101111111:	sigmoid_prime = 18'b001111101111111010;
		14'b11111110000000:	sigmoid_prime = 18'b001111110000001010;
		14'b11111110000001:	sigmoid_prime = 18'b001111110000011010;
		14'b11111110000010:	sigmoid_prime = 18'b001111110000101001;
		14'b11111110000011:	sigmoid_prime = 18'b001111110000111001;
		14'b11111110000100:	sigmoid_prime = 18'b001111110001001000;
		14'b11111110000101:	sigmoid_prime = 18'b001111110001010111;
		14'b11111110000110:	sigmoid_prime = 18'b001111110001100110;
		14'b11111110000111:	sigmoid_prime = 18'b001111110001110101;
		14'b11111110001000:	sigmoid_prime = 18'b001111110010000100;
		14'b11111110001001:	sigmoid_prime = 18'b001111110010010010;
		14'b11111110001010:	sigmoid_prime = 18'b001111110010100001;
		14'b11111110001011:	sigmoid_prime = 18'b001111110010101111;
		14'b11111110001100:	sigmoid_prime = 18'b001111110010111110;
		14'b11111110001101:	sigmoid_prime = 18'b001111110011001100;
		14'b11111110001110:	sigmoid_prime = 18'b001111110011011010;
		14'b11111110001111:	sigmoid_prime = 18'b001111110011101000;
		14'b11111110010000:	sigmoid_prime = 18'b001111110011110110;
		14'b11111110010001:	sigmoid_prime = 18'b001111110100000011;
		14'b11111110010010:	sigmoid_prime = 18'b001111110100010001;
		14'b11111110010011:	sigmoid_prime = 18'b001111110100011111;
		14'b11111110010100:	sigmoid_prime = 18'b001111110100101100;
		14'b11111110010101:	sigmoid_prime = 18'b001111110100111001;
		14'b11111110010110:	sigmoid_prime = 18'b001111110101000110;
		14'b11111110010111:	sigmoid_prime = 18'b001111110101010011;
		14'b11111110011000:	sigmoid_prime = 18'b001111110101100000;
		14'b11111110011001:	sigmoid_prime = 18'b001111110101101101;
		14'b11111110011010:	sigmoid_prime = 18'b001111110101111010;
		14'b11111110011011:	sigmoid_prime = 18'b001111110110000110;
		14'b11111110011100:	sigmoid_prime = 18'b001111110110010010;
		14'b11111110011101:	sigmoid_prime = 18'b001111110110011111;
		14'b11111110011110:	sigmoid_prime = 18'b001111110110101011;
		14'b11111110011111:	sigmoid_prime = 18'b001111110110110111;
		14'b11111110100000:	sigmoid_prime = 18'b001111110111000011;
		14'b11111110100001:	sigmoid_prime = 18'b001111110111001111;
		14'b11111110100010:	sigmoid_prime = 18'b001111110111011010;
		14'b11111110100011:	sigmoid_prime = 18'b001111110111100110;
		14'b11111110100100:	sigmoid_prime = 18'b001111110111110001;
		14'b11111110100101:	sigmoid_prime = 18'b001111110111111101;
		14'b11111110100110:	sigmoid_prime = 18'b001111111000001000;
		14'b11111110100111:	sigmoid_prime = 18'b001111111000010011;
		14'b11111110101000:	sigmoid_prime = 18'b001111111000011110;
		14'b11111110101001:	sigmoid_prime = 18'b001111111000101001;
		14'b11111110101010:	sigmoid_prime = 18'b001111111000110011;
		14'b11111110101011:	sigmoid_prime = 18'b001111111000111110;
		14'b11111110101100:	sigmoid_prime = 18'b001111111001001000;
		14'b11111110101101:	sigmoid_prime = 18'b001111111001010011;
		14'b11111110101110:	sigmoid_prime = 18'b001111111001011101;
		14'b11111110101111:	sigmoid_prime = 18'b001111111001100111;
		14'b11111110110000:	sigmoid_prime = 18'b001111111001110001;
		14'b11111110110001:	sigmoid_prime = 18'b001111111001111011;
		14'b11111110110010:	sigmoid_prime = 18'b001111111010000101;
		14'b11111110110011:	sigmoid_prime = 18'b001111111010001110;
		14'b11111110110100:	sigmoid_prime = 18'b001111111010011000;
		14'b11111110110101:	sigmoid_prime = 18'b001111111010100001;
		14'b11111110110110:	sigmoid_prime = 18'b001111111010101010;
		14'b11111110110111:	sigmoid_prime = 18'b001111111010110100;
		14'b11111110111000:	sigmoid_prime = 18'b001111111010111101;
		14'b11111110111001:	sigmoid_prime = 18'b001111111011000101;
		14'b11111110111010:	sigmoid_prime = 18'b001111111011001110;
		14'b11111110111011:	sigmoid_prime = 18'b001111111011010111;
		14'b11111110111100:	sigmoid_prime = 18'b001111111011011111;
		14'b11111110111101:	sigmoid_prime = 18'b001111111011101000;
		14'b11111110111110:	sigmoid_prime = 18'b001111111011110000;
		14'b11111110111111:	sigmoid_prime = 18'b001111111011111000;
		14'b11111111000000:	sigmoid_prime = 18'b001111111100000000;
		14'b11111111000001:	sigmoid_prime = 18'b001111111100001000;
		14'b11111111000010:	sigmoid_prime = 18'b001111111100010000;
		14'b11111111000011:	sigmoid_prime = 18'b001111111100010111;
		14'b11111111000100:	sigmoid_prime = 18'b001111111100011111;
		14'b11111111000101:	sigmoid_prime = 18'b001111111100100110;
		14'b11111111000110:	sigmoid_prime = 18'b001111111100101110;
		14'b11111111000111:	sigmoid_prime = 18'b001111111100110101;
		14'b11111111001000:	sigmoid_prime = 18'b001111111100111100;
		14'b11111111001001:	sigmoid_prime = 18'b001111111101000011;
		14'b11111111001010:	sigmoid_prime = 18'b001111111101001010;
		14'b11111111001011:	sigmoid_prime = 18'b001111111101010000;
		14'b11111111001100:	sigmoid_prime = 18'b001111111101010111;
		14'b11111111001101:	sigmoid_prime = 18'b001111111101011101;
		14'b11111111001110:	sigmoid_prime = 18'b001111111101100011;
		14'b11111111001111:	sigmoid_prime = 18'b001111111101101010;
		14'b11111111010000:	sigmoid_prime = 18'b001111111101110000;
		14'b11111111010001:	sigmoid_prime = 18'b001111111101110110;
		14'b11111111010010:	sigmoid_prime = 18'b001111111101111011;
		14'b11111111010011:	sigmoid_prime = 18'b001111111110000001;
		14'b11111111010100:	sigmoid_prime = 18'b001111111110000111;
		14'b11111111010101:	sigmoid_prime = 18'b001111111110001100;
		14'b11111111010110:	sigmoid_prime = 18'b001111111110010001;
		14'b11111111010111:	sigmoid_prime = 18'b001111111110010111;
		14'b11111111011000:	sigmoid_prime = 18'b001111111110011100;
		14'b11111111011001:	sigmoid_prime = 18'b001111111110100001;
		14'b11111111011010:	sigmoid_prime = 18'b001111111110100101;
		14'b11111111011011:	sigmoid_prime = 18'b001111111110101010;
		14'b11111111011100:	sigmoid_prime = 18'b001111111110101111;
		14'b11111111011101:	sigmoid_prime = 18'b001111111110110011;
		14'b11111111011110:	sigmoid_prime = 18'b001111111110110111;
		14'b11111111011111:	sigmoid_prime = 18'b001111111110111011;
		14'b11111111100000:	sigmoid_prime = 18'b001111111111000000;
		14'b11111111100001:	sigmoid_prime = 18'b001111111111000011;
		14'b11111111100010:	sigmoid_prime = 18'b001111111111000111;
		14'b11111111100011:	sigmoid_prime = 18'b001111111111001011;
		14'b11111111100100:	sigmoid_prime = 18'b001111111111001111;
		14'b11111111100101:	sigmoid_prime = 18'b001111111111010010;
		14'b11111111100110:	sigmoid_prime = 18'b001111111111010101;
		14'b11111111100111:	sigmoid_prime = 18'b001111111111011000;
		14'b11111111101000:	sigmoid_prime = 18'b001111111111011100;
		14'b11111111101001:	sigmoid_prime = 18'b001111111111011110;
		14'b11111111101010:	sigmoid_prime = 18'b001111111111100001;
		14'b11111111101011:	sigmoid_prime = 18'b001111111111100100;
		14'b11111111101100:	sigmoid_prime = 18'b001111111111100111;
		14'b11111111101101:	sigmoid_prime = 18'b001111111111101001;
		14'b11111111101110:	sigmoid_prime = 18'b001111111111101011;
		14'b11111111101111:	sigmoid_prime = 18'b001111111111101101;
		14'b11111111110000:	sigmoid_prime = 18'b001111111111110000;
		14'b11111111110001:	sigmoid_prime = 18'b001111111111110001;
		14'b11111111110010:	sigmoid_prime = 18'b001111111111110011;
		14'b11111111110011:	sigmoid_prime = 18'b001111111111110101;
		14'b11111111110100:	sigmoid_prime = 18'b001111111111110111;
		14'b11111111110101:	sigmoid_prime = 18'b001111111111111000;
		14'b11111111110110:	sigmoid_prime = 18'b001111111111111001;
		14'b11111111110111:	sigmoid_prime = 18'b001111111111111010;
		14'b11111111111000:	sigmoid_prime = 18'b001111111111111100;
		14'b11111111111001:	sigmoid_prime = 18'b001111111111111100;
		14'b11111111111010:	sigmoid_prime = 18'b001111111111111101;
		14'b11111111111011:	sigmoid_prime = 18'b001111111111111110;
		14'b11111111111100:	sigmoid_prime = 18'b001111111111111111;
		14'b11111111111101:	sigmoid_prime = 18'b001111111111111111;
		14'b11111111111110:	sigmoid_prime = 18'b001111111111111111;
		14'b11111111111111:	sigmoid_prime = 18'b001111111111111111;
		14'b00000000000000:	sigmoid_prime = 18'b010000000000000000;
		14'b00000000000001:	sigmoid_prime = 18'b001111111111111111;
		14'b00000000000010:	sigmoid_prime = 18'b001111111111111111;
		14'b00000000000011:	sigmoid_prime = 18'b001111111111111111;
		14'b00000000000100:	sigmoid_prime = 18'b001111111111111111;
		14'b00000000000101:	sigmoid_prime = 18'b001111111111111110;
		14'b00000000000110:	sigmoid_prime = 18'b001111111111111101;
		14'b00000000000111:	sigmoid_prime = 18'b001111111111111100;
		14'b00000000001000:	sigmoid_prime = 18'b001111111111111100;
		14'b00000000001001:	sigmoid_prime = 18'b001111111111111010;
		14'b00000000001010:	sigmoid_prime = 18'b001111111111111001;
		14'b00000000001011:	sigmoid_prime = 18'b001111111111111000;
		14'b00000000001100:	sigmoid_prime = 18'b001111111111110111;
		14'b00000000001101:	sigmoid_prime = 18'b001111111111110101;
		14'b00000000001110:	sigmoid_prime = 18'b001111111111110011;
		14'b00000000001111:	sigmoid_prime = 18'b001111111111110001;
		14'b00000000010000:	sigmoid_prime = 18'b001111111111110000;
		14'b00000000010001:	sigmoid_prime = 18'b001111111111101101;
		14'b00000000010010:	sigmoid_prime = 18'b001111111111101011;
		14'b00000000010011:	sigmoid_prime = 18'b001111111111101001;
		14'b00000000010100:	sigmoid_prime = 18'b001111111111100111;
		14'b00000000010101:	sigmoid_prime = 18'b001111111111100100;
		14'b00000000010110:	sigmoid_prime = 18'b001111111111100001;
		14'b00000000010111:	sigmoid_prime = 18'b001111111111011110;
		14'b00000000011000:	sigmoid_prime = 18'b001111111111011100;
		14'b00000000011001:	sigmoid_prime = 18'b001111111111011000;
		14'b00000000011010:	sigmoid_prime = 18'b001111111111010101;
		14'b00000000011011:	sigmoid_prime = 18'b001111111111010010;
		14'b00000000011100:	sigmoid_prime = 18'b001111111111001111;
		14'b00000000011101:	sigmoid_prime = 18'b001111111111001011;
		14'b00000000011110:	sigmoid_prime = 18'b001111111111000111;
		14'b00000000011111:	sigmoid_prime = 18'b001111111111000011;
		14'b00000000100000:	sigmoid_prime = 18'b001111111111000000;
		14'b00000000100001:	sigmoid_prime = 18'b001111111110111011;
		14'b00000000100010:	sigmoid_prime = 18'b001111111110110111;
		14'b00000000100011:	sigmoid_prime = 18'b001111111110110011;
		14'b00000000100100:	sigmoid_prime = 18'b001111111110101111;
		14'b00000000100101:	sigmoid_prime = 18'b001111111110101010;
		14'b00000000100110:	sigmoid_prime = 18'b001111111110100101;
		14'b00000000100111:	sigmoid_prime = 18'b001111111110100001;
		14'b00000000101000:	sigmoid_prime = 18'b001111111110011100;
		14'b00000000101001:	sigmoid_prime = 18'b001111111110010111;
		14'b00000000101010:	sigmoid_prime = 18'b001111111110010001;
		14'b00000000101011:	sigmoid_prime = 18'b001111111110001100;
		14'b00000000101100:	sigmoid_prime = 18'b001111111110000111;
		14'b00000000101101:	sigmoid_prime = 18'b001111111110000001;
		14'b00000000101110:	sigmoid_prime = 18'b001111111101111011;
		14'b00000000101111:	sigmoid_prime = 18'b001111111101110110;
		14'b00000000110000:	sigmoid_prime = 18'b001111111101110000;
		14'b00000000110001:	sigmoid_prime = 18'b001111111101101010;
		14'b00000000110010:	sigmoid_prime = 18'b001111111101100011;
		14'b00000000110011:	sigmoid_prime = 18'b001111111101011101;
		14'b00000000110100:	sigmoid_prime = 18'b001111111101010111;
		14'b00000000110101:	sigmoid_prime = 18'b001111111101010000;
		14'b00000000110110:	sigmoid_prime = 18'b001111111101001010;
		14'b00000000110111:	sigmoid_prime = 18'b001111111101000011;
		14'b00000000111000:	sigmoid_prime = 18'b001111111100111100;
		14'b00000000111001:	sigmoid_prime = 18'b001111111100110101;
		14'b00000000111010:	sigmoid_prime = 18'b001111111100101110;
		14'b00000000111011:	sigmoid_prime = 18'b001111111100100110;
		14'b00000000111100:	sigmoid_prime = 18'b001111111100011111;
		14'b00000000111101:	sigmoid_prime = 18'b001111111100010111;
		14'b00000000111110:	sigmoid_prime = 18'b001111111100010000;
		14'b00000000111111:	sigmoid_prime = 18'b001111111100001000;
		14'b00000001000000:	sigmoid_prime = 18'b001111111100000000;
		14'b00000001000001:	sigmoid_prime = 18'b001111111011111000;
		14'b00000001000010:	sigmoid_prime = 18'b001111111011110000;
		14'b00000001000011:	sigmoid_prime = 18'b001111111011101000;
		14'b00000001000100:	sigmoid_prime = 18'b001111111011011111;
		14'b00000001000101:	sigmoid_prime = 18'b001111111011010111;
		14'b00000001000110:	sigmoid_prime = 18'b001111111011001110;
		14'b00000001000111:	sigmoid_prime = 18'b001111111011000101;
		14'b00000001001000:	sigmoid_prime = 18'b001111111010111101;
		14'b00000001001001:	sigmoid_prime = 18'b001111111010110100;
		14'b00000001001010:	sigmoid_prime = 18'b001111111010101010;
		14'b00000001001011:	sigmoid_prime = 18'b001111111010100001;
		14'b00000001001100:	sigmoid_prime = 18'b001111111010011000;
		14'b00000001001101:	sigmoid_prime = 18'b001111111010001110;
		14'b00000001001110:	sigmoid_prime = 18'b001111111010000101;
		14'b00000001001111:	sigmoid_prime = 18'b001111111001111011;
		14'b00000001010000:	sigmoid_prime = 18'b001111111001110001;
		14'b00000001010001:	sigmoid_prime = 18'b001111111001100111;
		14'b00000001010010:	sigmoid_prime = 18'b001111111001011101;
		14'b00000001010011:	sigmoid_prime = 18'b001111111001010011;
		14'b00000001010100:	sigmoid_prime = 18'b001111111001001000;
		14'b00000001010101:	sigmoid_prime = 18'b001111111000111110;
		14'b00000001010110:	sigmoid_prime = 18'b001111111000110011;
		14'b00000001010111:	sigmoid_prime = 18'b001111111000101001;
		14'b00000001011000:	sigmoid_prime = 18'b001111111000011110;
		14'b00000001011001:	sigmoid_prime = 18'b001111111000010011;
		14'b00000001011010:	sigmoid_prime = 18'b001111111000001000;
		14'b00000001011011:	sigmoid_prime = 18'b001111110111111101;
		14'b00000001011100:	sigmoid_prime = 18'b001111110111110001;
		14'b00000001011101:	sigmoid_prime = 18'b001111110111100110;
		14'b00000001011110:	sigmoid_prime = 18'b001111110111011010;
		14'b00000001011111:	sigmoid_prime = 18'b001111110111001111;
		14'b00000001100000:	sigmoid_prime = 18'b001111110111000011;
		14'b00000001100001:	sigmoid_prime = 18'b001111110110110111;
		14'b00000001100010:	sigmoid_prime = 18'b001111110110101011;
		14'b00000001100011:	sigmoid_prime = 18'b001111110110011111;
		14'b00000001100100:	sigmoid_prime = 18'b001111110110010010;
		14'b00000001100101:	sigmoid_prime = 18'b001111110110000110;
		14'b00000001100110:	sigmoid_prime = 18'b001111110101111010;
		14'b00000001100111:	sigmoid_prime = 18'b001111110101101101;
		14'b00000001101000:	sigmoid_prime = 18'b001111110101100000;
		14'b00000001101001:	sigmoid_prime = 18'b001111110101010011;
		14'b00000001101010:	sigmoid_prime = 18'b001111110101000110;
		14'b00000001101011:	sigmoid_prime = 18'b001111110100111001;
		14'b00000001101100:	sigmoid_prime = 18'b001111110100101100;
		14'b00000001101101:	sigmoid_prime = 18'b001111110100011111;
		14'b00000001101110:	sigmoid_prime = 18'b001111110100010001;
		14'b00000001101111:	sigmoid_prime = 18'b001111110100000011;
		14'b00000001110000:	sigmoid_prime = 18'b001111110011110110;
		14'b00000001110001:	sigmoid_prime = 18'b001111110011101000;
		14'b00000001110010:	sigmoid_prime = 18'b001111110011011010;
		14'b00000001110011:	sigmoid_prime = 18'b001111110011001100;
		14'b00000001110100:	sigmoid_prime = 18'b001111110010111110;
		14'b00000001110101:	sigmoid_prime = 18'b001111110010101111;
		14'b00000001110110:	sigmoid_prime = 18'b001111110010100001;
		14'b00000001110111:	sigmoid_prime = 18'b001111110010010010;
		14'b00000001111000:	sigmoid_prime = 18'b001111110010000100;
		14'b00000001111001:	sigmoid_prime = 18'b001111110001110101;
		14'b00000001111010:	sigmoid_prime = 18'b001111110001100110;
		14'b00000001111011:	sigmoid_prime = 18'b001111110001010111;
		14'b00000001111100:	sigmoid_prime = 18'b001111110001001000;
		14'b00000001111101:	sigmoid_prime = 18'b001111110000111001;
		14'b00000001111110:	sigmoid_prime = 18'b001111110000101001;
		14'b00000001111111:	sigmoid_prime = 18'b001111110000011010;
		14'b00000010000000:	sigmoid_prime = 18'b001111110000001010;
		14'b00000010000001:	sigmoid_prime = 18'b001111101111111010;
		14'b00000010000010:	sigmoid_prime = 18'b001111101111101010;
		14'b00000010000011:	sigmoid_prime = 18'b001111101111011011;
		14'b00000010000100:	sigmoid_prime = 18'b001111101111001010;
		14'b00000010000101:	sigmoid_prime = 18'b001111101110111010;
		14'b00000010000110:	sigmoid_prime = 18'b001111101110101010;
		14'b00000010000111:	sigmoid_prime = 18'b001111101110011010;
		14'b00000010001000:	sigmoid_prime = 18'b001111101110001001;
		14'b00000010001001:	sigmoid_prime = 18'b001111101101111000;
		14'b00000010001010:	sigmoid_prime = 18'b001111101101101000;
		14'b00000010001011:	sigmoid_prime = 18'b001111101101010111;
		14'b00000010001100:	sigmoid_prime = 18'b001111101101000110;
		14'b00000010001101:	sigmoid_prime = 18'b001111101100110100;
		14'b00000010001110:	sigmoid_prime = 18'b001111101100100011;
		14'b00000010001111:	sigmoid_prime = 18'b001111101100010010;
		14'b00000010010000:	sigmoid_prime = 18'b001111101100000000;
		14'b00000010010001:	sigmoid_prime = 18'b001111101011101111;
		14'b00000010010010:	sigmoid_prime = 18'b001111101011011101;
		14'b00000010010011:	sigmoid_prime = 18'b001111101011001011;
		14'b00000010010100:	sigmoid_prime = 18'b001111101010111001;
		14'b00000010010101:	sigmoid_prime = 18'b001111101010100111;
		14'b00000010010110:	sigmoid_prime = 18'b001111101010010101;
		14'b00000010010111:	sigmoid_prime = 18'b001111101010000011;
		14'b00000010011000:	sigmoid_prime = 18'b001111101001110000;
		14'b00000010011001:	sigmoid_prime = 18'b001111101001011110;
		14'b00000010011010:	sigmoid_prime = 18'b001111101001001011;
		14'b00000010011011:	sigmoid_prime = 18'b001111101000111001;
		14'b00000010011100:	sigmoid_prime = 18'b001111101000100110;
		14'b00000010011101:	sigmoid_prime = 18'b001111101000010011;
		14'b00000010011110:	sigmoid_prime = 18'b001111101000000000;
		14'b00000010011111:	sigmoid_prime = 18'b001111100111101100;
		14'b00000010100000:	sigmoid_prime = 18'b001111100111011001;
		14'b00000010100001:	sigmoid_prime = 18'b001111100111000110;
		14'b00000010100010:	sigmoid_prime = 18'b001111100110110010;
		14'b00000010100011:	sigmoid_prime = 18'b001111100110011111;
		14'b00000010100100:	sigmoid_prime = 18'b001111100110001011;
		14'b00000010100101:	sigmoid_prime = 18'b001111100101110111;
		14'b00000010100110:	sigmoid_prime = 18'b001111100101100011;
		14'b00000010100111:	sigmoid_prime = 18'b001111100101001111;
		14'b00000010101000:	sigmoid_prime = 18'b001111100100111011;
		14'b00000010101001:	sigmoid_prime = 18'b001111100100100110;
		14'b00000010101010:	sigmoid_prime = 18'b001111100100010010;
		14'b00000010101011:	sigmoid_prime = 18'b001111100011111101;
		14'b00000010101100:	sigmoid_prime = 18'b001111100011101001;
		14'b00000010101101:	sigmoid_prime = 18'b001111100011010100;
		14'b00000010101110:	sigmoid_prime = 18'b001111100010111111;
		14'b00000010101111:	sigmoid_prime = 18'b001111100010101010;
		14'b00000010110000:	sigmoid_prime = 18'b001111100010010101;
		14'b00000010110001:	sigmoid_prime = 18'b001111100010000000;
		14'b00000010110010:	sigmoid_prime = 18'b001111100001101010;
		14'b00000010110011:	sigmoid_prime = 18'b001111100001010101;
		14'b00000010110100:	sigmoid_prime = 18'b001111100000111111;
		14'b00000010110101:	sigmoid_prime = 18'b001111100000101010;
		14'b00000010110110:	sigmoid_prime = 18'b001111100000010100;
		14'b00000010110111:	sigmoid_prime = 18'b001111011111111110;
		14'b00000010111000:	sigmoid_prime = 18'b001111011111101000;
		14'b00000010111001:	sigmoid_prime = 18'b001111011111010010;
		14'b00000010111010:	sigmoid_prime = 18'b001111011110111100;
		14'b00000010111011:	sigmoid_prime = 18'b001111011110100110;
		14'b00000010111100:	sigmoid_prime = 18'b001111011110001111;
		14'b00000010111101:	sigmoid_prime = 18'b001111011101111001;
		14'b00000010111110:	sigmoid_prime = 18'b001111011101100010;
		14'b00000010111111:	sigmoid_prime = 18'b001111011101001011;
		14'b00000011000000:	sigmoid_prime = 18'b001111011100110100;
		14'b00000011000001:	sigmoid_prime = 18'b001111011100011101;
		14'b00000011000010:	sigmoid_prime = 18'b001111011100000110;
		14'b00000011000011:	sigmoid_prime = 18'b001111011011101111;
		14'b00000011000100:	sigmoid_prime = 18'b001111011011011000;
		14'b00000011000101:	sigmoid_prime = 18'b001111011011000001;
		14'b00000011000110:	sigmoid_prime = 18'b001111011010101001;
		14'b00000011000111:	sigmoid_prime = 18'b001111011010010001;
		14'b00000011001000:	sigmoid_prime = 18'b001111011001111010;
		14'b00000011001001:	sigmoid_prime = 18'b001111011001100010;
		14'b00000011001010:	sigmoid_prime = 18'b001111011001001010;
		14'b00000011001011:	sigmoid_prime = 18'b001111011000110010;
		14'b00000011001100:	sigmoid_prime = 18'b001111011000011010;
		14'b00000011001101:	sigmoid_prime = 18'b001111011000000010;
		14'b00000011001110:	sigmoid_prime = 18'b001111010111101001;
		14'b00000011001111:	sigmoid_prime = 18'b001111010111010001;
		14'b00000011010000:	sigmoid_prime = 18'b001111010110111000;
		14'b00000011010001:	sigmoid_prime = 18'b001111010110100000;
		14'b00000011010010:	sigmoid_prime = 18'b001111010110000111;
		14'b00000011010011:	sigmoid_prime = 18'b001111010101101110;
		14'b00000011010100:	sigmoid_prime = 18'b001111010101010101;
		14'b00000011010101:	sigmoid_prime = 18'b001111010100111100;
		14'b00000011010110:	sigmoid_prime = 18'b001111010100100011;
		14'b00000011010111:	sigmoid_prime = 18'b001111010100001001;
		14'b00000011011000:	sigmoid_prime = 18'b001111010011110000;
		14'b00000011011001:	sigmoid_prime = 18'b001111010011010110;
		14'b00000011011010:	sigmoid_prime = 18'b001111010010111101;
		14'b00000011011011:	sigmoid_prime = 18'b001111010010100011;
		14'b00000011011100:	sigmoid_prime = 18'b001111010010001001;
		14'b00000011011101:	sigmoid_prime = 18'b001111010001101111;
		14'b00000011011110:	sigmoid_prime = 18'b001111010001010101;
		14'b00000011011111:	sigmoid_prime = 18'b001111010000111011;
		14'b00000011100000:	sigmoid_prime = 18'b001111010000100001;
		14'b00000011100001:	sigmoid_prime = 18'b001111010000000111;
		14'b00000011100010:	sigmoid_prime = 18'b001111001111101100;
		14'b00000011100011:	sigmoid_prime = 18'b001111001111010010;
		14'b00000011100100:	sigmoid_prime = 18'b001111001110110111;
		14'b00000011100101:	sigmoid_prime = 18'b001111001110011100;
		14'b00000011100110:	sigmoid_prime = 18'b001111001110000001;
		14'b00000011100111:	sigmoid_prime = 18'b001111001101100110;
		14'b00000011101000:	sigmoid_prime = 18'b001111001101001011;
		14'b00000011101001:	sigmoid_prime = 18'b001111001100110000;
		14'b00000011101010:	sigmoid_prime = 18'b001111001100010101;
		14'b00000011101011:	sigmoid_prime = 18'b001111001011111010;
		14'b00000011101100:	sigmoid_prime = 18'b001111001011011110;
		14'b00000011101101:	sigmoid_prime = 18'b001111001011000011;
		14'b00000011101110:	sigmoid_prime = 18'b001111001010100111;
		14'b00000011101111:	sigmoid_prime = 18'b001111001010001011;
		14'b00000011110000:	sigmoid_prime = 18'b001111001001101111;
		14'b00000011110001:	sigmoid_prime = 18'b001111001001010011;
		14'b00000011110010:	sigmoid_prime = 18'b001111001000110111;
		14'b00000011110011:	sigmoid_prime = 18'b001111001000011011;
		14'b00000011110100:	sigmoid_prime = 18'b001111000111111111;
		14'b00000011110101:	sigmoid_prime = 18'b001111000111100011;
		14'b00000011110110:	sigmoid_prime = 18'b001111000111000110;
		14'b00000011110111:	sigmoid_prime = 18'b001111000110101010;
		14'b00000011111000:	sigmoid_prime = 18'b001111000110001101;
		14'b00000011111001:	sigmoid_prime = 18'b001111000101110000;
		14'b00000011111010:	sigmoid_prime = 18'b001111000101010011;
		14'b00000011111011:	sigmoid_prime = 18'b001111000100110110;
		14'b00000011111100:	sigmoid_prime = 18'b001111000100011001;
		14'b00000011111101:	sigmoid_prime = 18'b001111000011111100;
		14'b00000011111110:	sigmoid_prime = 18'b001111000011011111;
		14'b00000011111111:	sigmoid_prime = 18'b001111000011000010;
		14'b00000100000000:	sigmoid_prime = 18'b001111000010100100;
		14'b00000100000001:	sigmoid_prime = 18'b001111000010000111;
		14'b00000100000010:	sigmoid_prime = 18'b001111000001101001;
		14'b00000100000011:	sigmoid_prime = 18'b001111000001001011;
		14'b00000100000100:	sigmoid_prime = 18'b001111000000101110;
		14'b00000100000101:	sigmoid_prime = 18'b001111000000010000;
		14'b00000100000110:	sigmoid_prime = 18'b001110111111110010;
		14'b00000100000111:	sigmoid_prime = 18'b001110111111010100;
		14'b00000100001000:	sigmoid_prime = 18'b001110111110110101;
		14'b00000100001001:	sigmoid_prime = 18'b001110111110010111;
		14'b00000100001010:	sigmoid_prime = 18'b001110111101111001;
		14'b00000100001011:	sigmoid_prime = 18'b001110111101011010;
		14'b00000100001100:	sigmoid_prime = 18'b001110111100111100;
		14'b00000100001101:	sigmoid_prime = 18'b001110111100011101;
		14'b00000100001110:	sigmoid_prime = 18'b001110111011111110;
		14'b00000100001111:	sigmoid_prime = 18'b001110111011100000;
		14'b00000100010000:	sigmoid_prime = 18'b001110111011000001;
		14'b00000100010001:	sigmoid_prime = 18'b001110111010100010;
		14'b00000100010010:	sigmoid_prime = 18'b001110111010000010;
		14'b00000100010011:	sigmoid_prime = 18'b001110111001100011;
		14'b00000100010100:	sigmoid_prime = 18'b001110111001000100;
		14'b00000100010101:	sigmoid_prime = 18'b001110111000100101;
		14'b00000100010110:	sigmoid_prime = 18'b001110111000000101;
		14'b00000100010111:	sigmoid_prime = 18'b001110110111100101;
		14'b00000100011000:	sigmoid_prime = 18'b001110110111000110;
		14'b00000100011001:	sigmoid_prime = 18'b001110110110100110;
		14'b00000100011010:	sigmoid_prime = 18'b001110110110000110;
		14'b00000100011011:	sigmoid_prime = 18'b001110110101100110;
		14'b00000100011100:	sigmoid_prime = 18'b001110110101000110;
		14'b00000100011101:	sigmoid_prime = 18'b001110110100100110;
		14'b00000100011110:	sigmoid_prime = 18'b001110110100000110;
		14'b00000100011111:	sigmoid_prime = 18'b001110110011100110;
		14'b00000100100000:	sigmoid_prime = 18'b001110110011000101;
		14'b00000100100001:	sigmoid_prime = 18'b001110110010100101;
		14'b00000100100010:	sigmoid_prime = 18'b001110110010000100;
		14'b00000100100011:	sigmoid_prime = 18'b001110110001100011;
		14'b00000100100100:	sigmoid_prime = 18'b001110110001000011;
		14'b00000100100101:	sigmoid_prime = 18'b001110110000100010;
		14'b00000100100110:	sigmoid_prime = 18'b001110110000000001;
		14'b00000100100111:	sigmoid_prime = 18'b001110101111100000;
		14'b00000100101000:	sigmoid_prime = 18'b001110101110111111;
		14'b00000100101001:	sigmoid_prime = 18'b001110101110011110;
		14'b00000100101010:	sigmoid_prime = 18'b001110101101111100;
		14'b00000100101011:	sigmoid_prime = 18'b001110101101011011;
		14'b00000100101100:	sigmoid_prime = 18'b001110101100111001;
		14'b00000100101101:	sigmoid_prime = 18'b001110101100011000;
		14'b00000100101110:	sigmoid_prime = 18'b001110101011110110;
		14'b00000100101111:	sigmoid_prime = 18'b001110101011010100;
		14'b00000100110000:	sigmoid_prime = 18'b001110101010110011;
		14'b00000100110001:	sigmoid_prime = 18'b001110101010010001;
		14'b00000100110010:	sigmoid_prime = 18'b001110101001101111;
		14'b00000100110011:	sigmoid_prime = 18'b001110101001001101;
		14'b00000100110100:	sigmoid_prime = 18'b001110101000101011;
		14'b00000100110101:	sigmoid_prime = 18'b001110101000001000;
		14'b00000100110110:	sigmoid_prime = 18'b001110100111100110;
		14'b00000100110111:	sigmoid_prime = 18'b001110100111000100;
		14'b00000100111000:	sigmoid_prime = 18'b001110100110100001;
		14'b00000100111001:	sigmoid_prime = 18'b001110100101111111;
		14'b00000100111010:	sigmoid_prime = 18'b001110100101011100;
		14'b00000100111011:	sigmoid_prime = 18'b001110100100111001;
		14'b00000100111100:	sigmoid_prime = 18'b001110100100010110;
		14'b00000100111101:	sigmoid_prime = 18'b001110100011110011;
		14'b00000100111110:	sigmoid_prime = 18'b001110100011010000;
		14'b00000100111111:	sigmoid_prime = 18'b001110100010101101;
		14'b00000101000000:	sigmoid_prime = 18'b001110100010001010;
		14'b00000101000001:	sigmoid_prime = 18'b001110100001100111;
		14'b00000101000010:	sigmoid_prime = 18'b001110100001000100;
		14'b00000101000011:	sigmoid_prime = 18'b001110100000100000;
		14'b00000101000100:	sigmoid_prime = 18'b001110011111111101;
		14'b00000101000101:	sigmoid_prime = 18'b001110011111011001;
		14'b00000101000110:	sigmoid_prime = 18'b001110011110110110;
		14'b00000101000111:	sigmoid_prime = 18'b001110011110010010;
		14'b00000101001000:	sigmoid_prime = 18'b001110011101101110;
		14'b00000101001001:	sigmoid_prime = 18'b001110011101001010;
		14'b00000101001010:	sigmoid_prime = 18'b001110011100100110;
		14'b00000101001011:	sigmoid_prime = 18'b001110011100000010;
		14'b00000101001100:	sigmoid_prime = 18'b001110011011011110;
		14'b00000101001101:	sigmoid_prime = 18'b001110011010111010;
		14'b00000101001110:	sigmoid_prime = 18'b001110011010010110;
		14'b00000101001111:	sigmoid_prime = 18'b001110011001110001;
		14'b00000101010000:	sigmoid_prime = 18'b001110011001001101;
		14'b00000101010001:	sigmoid_prime = 18'b001110011000101000;
		14'b00000101010010:	sigmoid_prime = 18'b001110011000000100;
		14'b00000101010011:	sigmoid_prime = 18'b001110010111011111;
		14'b00000101010100:	sigmoid_prime = 18'b001110010110111010;
		14'b00000101010101:	sigmoid_prime = 18'b001110010110010101;
		14'b00000101010110:	sigmoid_prime = 18'b001110010101110000;
		14'b00000101010111:	sigmoid_prime = 18'b001110010101001011;
		14'b00000101011000:	sigmoid_prime = 18'b001110010100100110;
		14'b00000101011001:	sigmoid_prime = 18'b001110010100000001;
		14'b00000101011010:	sigmoid_prime = 18'b001110010011011100;
		14'b00000101011011:	sigmoid_prime = 18'b001110010010110111;
		14'b00000101011100:	sigmoid_prime = 18'b001110010010010001;
		14'b00000101011101:	sigmoid_prime = 18'b001110010001101100;
		14'b00000101011110:	sigmoid_prime = 18'b001110010001000110;
		14'b00000101011111:	sigmoid_prime = 18'b001110010000100001;
		14'b00000101100000:	sigmoid_prime = 18'b001110001111111011;
		14'b00000101100001:	sigmoid_prime = 18'b001110001111010101;
		14'b00000101100010:	sigmoid_prime = 18'b001110001110101111;
		14'b00000101100011:	sigmoid_prime = 18'b001110001110001010;
		14'b00000101100100:	sigmoid_prime = 18'b001110001101100100;
		14'b00000101100101:	sigmoid_prime = 18'b001110001100111110;
		14'b00000101100110:	sigmoid_prime = 18'b001110001100010111;
		14'b00000101100111:	sigmoid_prime = 18'b001110001011110001;
		14'b00000101101000:	sigmoid_prime = 18'b001110001011001011;
		14'b00000101101001:	sigmoid_prime = 18'b001110001010100101;
		14'b00000101101010:	sigmoid_prime = 18'b001110001001111110;
		14'b00000101101011:	sigmoid_prime = 18'b001110001001011000;
		14'b00000101101100:	sigmoid_prime = 18'b001110001000110001;
		14'b00000101101101:	sigmoid_prime = 18'b001110001000001011;
		14'b00000101101110:	sigmoid_prime = 18'b001110000111100100;
		14'b00000101101111:	sigmoid_prime = 18'b001110000110111101;
		14'b00000101110000:	sigmoid_prime = 18'b001110000110010110;
		14'b00000101110001:	sigmoid_prime = 18'b001110000101101111;
		14'b00000101110010:	sigmoid_prime = 18'b001110000101001000;
		14'b00000101110011:	sigmoid_prime = 18'b001110000100100001;
		14'b00000101110100:	sigmoid_prime = 18'b001110000011111010;
		14'b00000101110101:	sigmoid_prime = 18'b001110000011010011;
		14'b00000101110110:	sigmoid_prime = 18'b001110000010101100;
		14'b00000101110111:	sigmoid_prime = 18'b001110000010000100;
		14'b00000101111000:	sigmoid_prime = 18'b001110000001011101;
		14'b00000101111001:	sigmoid_prime = 18'b001110000000110110;
		14'b00000101111010:	sigmoid_prime = 18'b001110000000001110;
		14'b00000101111011:	sigmoid_prime = 18'b001101111111100110;
		14'b00000101111100:	sigmoid_prime = 18'b001101111110111111;
		14'b00000101111101:	sigmoid_prime = 18'b001101111110010111;
		14'b00000101111110:	sigmoid_prime = 18'b001101111101101111;
		14'b00000101111111:	sigmoid_prime = 18'b001101111101000111;
		14'b00000110000000:	sigmoid_prime = 18'b001101111100011111;
		14'b00000110000001:	sigmoid_prime = 18'b001101111011110111;
		14'b00000110000010:	sigmoid_prime = 18'b001101111011001111;
		14'b00000110000011:	sigmoid_prime = 18'b001101111010100111;
		14'b00000110000100:	sigmoid_prime = 18'b001101111001111111;
		14'b00000110000101:	sigmoid_prime = 18'b001101111001010111;
		14'b00000110000110:	sigmoid_prime = 18'b001101111000101110;
		14'b00000110000111:	sigmoid_prime = 18'b001101111000000110;
		14'b00000110001000:	sigmoid_prime = 18'b001101110111011101;
		14'b00000110001001:	sigmoid_prime = 18'b001101110110110101;
		14'b00000110001010:	sigmoid_prime = 18'b001101110110001100;
		14'b00000110001011:	sigmoid_prime = 18'b001101110101100100;
		14'b00000110001100:	sigmoid_prime = 18'b001101110100111011;
		14'b00000110001101:	sigmoid_prime = 18'b001101110100010010;
		14'b00000110001110:	sigmoid_prime = 18'b001101110011101001;
		14'b00000110001111:	sigmoid_prime = 18'b001101110011000000;
		14'b00000110010000:	sigmoid_prime = 18'b001101110010010111;
		14'b00000110010001:	sigmoid_prime = 18'b001101110001101110;
		14'b00000110010010:	sigmoid_prime = 18'b001101110001000101;
		14'b00000110010011:	sigmoid_prime = 18'b001101110000011100;
		14'b00000110010100:	sigmoid_prime = 18'b001101101111110011;
		14'b00000110010101:	sigmoid_prime = 18'b001101101111001001;
		14'b00000110010110:	sigmoid_prime = 18'b001101101110100000;
		14'b00000110010111:	sigmoid_prime = 18'b001101101101110111;
		14'b00000110011000:	sigmoid_prime = 18'b001101101101001101;
		14'b00000110011001:	sigmoid_prime = 18'b001101101100100100;
		14'b00000110011010:	sigmoid_prime = 18'b001101101011111010;
		14'b00000110011011:	sigmoid_prime = 18'b001101101011010000;
		14'b00000110011100:	sigmoid_prime = 18'b001101101010100111;
		14'b00000110011101:	sigmoid_prime = 18'b001101101001111101;
		14'b00000110011110:	sigmoid_prime = 18'b001101101001010011;
		14'b00000110011111:	sigmoid_prime = 18'b001101101000101001;
		14'b00000110100000:	sigmoid_prime = 18'b001101100111111111;
		14'b00000110100001:	sigmoid_prime = 18'b001101100111010101;
		14'b00000110100010:	sigmoid_prime = 18'b001101100110101011;
		14'b00000110100011:	sigmoid_prime = 18'b001101100110000001;
		14'b00000110100100:	sigmoid_prime = 18'b001101100101010111;
		14'b00000110100101:	sigmoid_prime = 18'b001101100100101100;
		14'b00000110100110:	sigmoid_prime = 18'b001101100100000010;
		14'b00000110100111:	sigmoid_prime = 18'b001101100011011000;
		14'b00000110101000:	sigmoid_prime = 18'b001101100010101101;
		14'b00000110101001:	sigmoid_prime = 18'b001101100010000011;
		14'b00000110101010:	sigmoid_prime = 18'b001101100001011000;
		14'b00000110101011:	sigmoid_prime = 18'b001101100000101110;
		14'b00000110101100:	sigmoid_prime = 18'b001101100000000011;
		14'b00000110101101:	sigmoid_prime = 18'b001101011111011000;
		14'b00000110101110:	sigmoid_prime = 18'b001101011110101101;
		14'b00000110101111:	sigmoid_prime = 18'b001101011110000011;
		14'b00000110110000:	sigmoid_prime = 18'b001101011101011000;
		14'b00000110110001:	sigmoid_prime = 18'b001101011100101101;
		14'b00000110110010:	sigmoid_prime = 18'b001101011100000010;
		14'b00000110110011:	sigmoid_prime = 18'b001101011011010111;
		14'b00000110110100:	sigmoid_prime = 18'b001101011010101100;
		14'b00000110110101:	sigmoid_prime = 18'b001101011010000001;
		14'b00000110110110:	sigmoid_prime = 18'b001101011001010101;
		14'b00000110110111:	sigmoid_prime = 18'b001101011000101010;
		14'b00000110111000:	sigmoid_prime = 18'b001101010111111111;
		14'b00000110111001:	sigmoid_prime = 18'b001101010111010011;
		14'b00000110111010:	sigmoid_prime = 18'b001101010110101000;
		14'b00000110111011:	sigmoid_prime = 18'b001101010101111101;
		14'b00000110111100:	sigmoid_prime = 18'b001101010101010001;
		14'b00000110111101:	sigmoid_prime = 18'b001101010100100101;
		14'b00000110111110:	sigmoid_prime = 18'b001101010011111010;
		14'b00000110111111:	sigmoid_prime = 18'b001101010011001110;
		14'b00000111000000:	sigmoid_prime = 18'b001101010010100010;
		14'b00000111000001:	sigmoid_prime = 18'b001101010001110111;
		14'b00000111000010:	sigmoid_prime = 18'b001101010001001011;
		14'b00000111000011:	sigmoid_prime = 18'b001101010000011111;
		14'b00000111000100:	sigmoid_prime = 18'b001101001111110011;
		14'b00000111000101:	sigmoid_prime = 18'b001101001111000111;
		14'b00000111000110:	sigmoid_prime = 18'b001101001110011011;
		14'b00000111000111:	sigmoid_prime = 18'b001101001101101111;
		14'b00000111001000:	sigmoid_prime = 18'b001101001101000011;
		14'b00000111001001:	sigmoid_prime = 18'b001101001100010111;
		14'b00000111001010:	sigmoid_prime = 18'b001101001011101010;
		14'b00000111001011:	sigmoid_prime = 18'b001101001010111110;
		14'b00000111001100:	sigmoid_prime = 18'b001101001010010010;
		14'b00000111001101:	sigmoid_prime = 18'b001101001001100101;
		14'b00000111001110:	sigmoid_prime = 18'b001101001000111001;
		14'b00000111001111:	sigmoid_prime = 18'b001101001000001100;
		14'b00000111010000:	sigmoid_prime = 18'b001101000111100000;
		14'b00000111010001:	sigmoid_prime = 18'b001101000110110011;
		14'b00000111010010:	sigmoid_prime = 18'b001101000110000111;
		14'b00000111010011:	sigmoid_prime = 18'b001101000101011010;
		14'b00000111010100:	sigmoid_prime = 18'b001101000100101101;
		14'b00000111010101:	sigmoid_prime = 18'b001101000100000001;
		14'b00000111010110:	sigmoid_prime = 18'b001101000011010100;
		14'b00000111010111:	sigmoid_prime = 18'b001101000010100111;
		14'b00000111011000:	sigmoid_prime = 18'b001101000001111010;
		14'b00000111011001:	sigmoid_prime = 18'b001101000001001101;
		14'b00000111011010:	sigmoid_prime = 18'b001101000000100000;
		14'b00000111011011:	sigmoid_prime = 18'b001100111111110011;
		14'b00000111011100:	sigmoid_prime = 18'b001100111111000110;
		14'b00000111011101:	sigmoid_prime = 18'b001100111110011001;
		14'b00000111011110:	sigmoid_prime = 18'b001100111101101100;
		14'b00000111011111:	sigmoid_prime = 18'b001100111100111111;
		14'b00000111100000:	sigmoid_prime = 18'b001100111100010001;
		14'b00000111100001:	sigmoid_prime = 18'b001100111011100100;
		14'b00000111100010:	sigmoid_prime = 18'b001100111010110111;
		14'b00000111100011:	sigmoid_prime = 18'b001100111010001001;
		14'b00000111100100:	sigmoid_prime = 18'b001100111001011100;
		14'b00000111100101:	sigmoid_prime = 18'b001100111000101110;
		14'b00000111100110:	sigmoid_prime = 18'b001100111000000001;
		14'b00000111100111:	sigmoid_prime = 18'b001100110111010011;
		14'b00000111101000:	sigmoid_prime = 18'b001100110110100110;
		14'b00000111101001:	sigmoid_prime = 18'b001100110101111000;
		14'b00000111101010:	sigmoid_prime = 18'b001100110101001011;
		14'b00000111101011:	sigmoid_prime = 18'b001100110100011101;
		14'b00000111101100:	sigmoid_prime = 18'b001100110011101111;
		14'b00000111101101:	sigmoid_prime = 18'b001100110011000001;
		14'b00000111101110:	sigmoid_prime = 18'b001100110010010100;
		14'b00000111101111:	sigmoid_prime = 18'b001100110001100110;
		14'b00000111110000:	sigmoid_prime = 18'b001100110000111000;
		14'b00000111110001:	sigmoid_prime = 18'b001100110000001010;
		14'b00000111110010:	sigmoid_prime = 18'b001100101111011100;
		14'b00000111110011:	sigmoid_prime = 18'b001100101110101110;
		14'b00000111110100:	sigmoid_prime = 18'b001100101110000000;
		14'b00000111110101:	sigmoid_prime = 18'b001100101101010010;
		14'b00000111110110:	sigmoid_prime = 18'b001100101100100100;
		14'b00000111110111:	sigmoid_prime = 18'b001100101011110101;
		14'b00000111111000:	sigmoid_prime = 18'b001100101011000111;
		14'b00000111111001:	sigmoid_prime = 18'b001100101010011001;
		14'b00000111111010:	sigmoid_prime = 18'b001100101001101011;
		14'b00000111111011:	sigmoid_prime = 18'b001100101000111100;
		14'b00000111111100:	sigmoid_prime = 18'b001100101000001110;
		14'b00000111111101:	sigmoid_prime = 18'b001100100111100000;
		14'b00000111111110:	sigmoid_prime = 18'b001100100110110001;
		14'b00000111111111:	sigmoid_prime = 18'b001100100110000011;
		14'b00001000000000:	sigmoid_prime = 18'b001100100101010100;
		14'b00001000000001:	sigmoid_prime = 18'b001100100100100110;
		14'b00001000000010:	sigmoid_prime = 18'b001100100011110111;
		14'b00001000000011:	sigmoid_prime = 18'b001100100011001000;
		14'b00001000000100:	sigmoid_prime = 18'b001100100010011010;
		14'b00001000000101:	sigmoid_prime = 18'b001100100001101011;
		14'b00001000000110:	sigmoid_prime = 18'b001100100000111100;
		14'b00001000000111:	sigmoid_prime = 18'b001100100000001110;
		14'b00001000001000:	sigmoid_prime = 18'b001100011111011111;
		14'b00001000001001:	sigmoid_prime = 18'b001100011110110000;
		14'b00001000001010:	sigmoid_prime = 18'b001100011110000001;
		14'b00001000001011:	sigmoid_prime = 18'b001100011101010010;
		14'b00001000001100:	sigmoid_prime = 18'b001100011100100011;
		14'b00001000001101:	sigmoid_prime = 18'b001100011011110100;
		14'b00001000001110:	sigmoid_prime = 18'b001100011011000110;
		14'b00001000001111:	sigmoid_prime = 18'b001100011010010111;
		14'b00001000010000:	sigmoid_prime = 18'b001100011001100111;
		14'b00001000010001:	sigmoid_prime = 18'b001100011000111000;
		14'b00001000010010:	sigmoid_prime = 18'b001100011000001001;
		14'b00001000010011:	sigmoid_prime = 18'b001100010111011010;
		14'b00001000010100:	sigmoid_prime = 18'b001100010110101011;
		14'b00001000010101:	sigmoid_prime = 18'b001100010101111100;
		14'b00001000010110:	sigmoid_prime = 18'b001100010101001101;
		14'b00001000010111:	sigmoid_prime = 18'b001100010100011101;
		14'b00001000011000:	sigmoid_prime = 18'b001100010011101110;
		14'b00001000011001:	sigmoid_prime = 18'b001100010010111111;
		14'b00001000011010:	sigmoid_prime = 18'b001100010010001111;
		14'b00001000011011:	sigmoid_prime = 18'b001100010001100000;
		14'b00001000011100:	sigmoid_prime = 18'b001100010000110001;
		14'b00001000011101:	sigmoid_prime = 18'b001100010000000001;
		14'b00001000011110:	sigmoid_prime = 18'b001100001111010010;
		14'b00001000011111:	sigmoid_prime = 18'b001100001110100010;
		14'b00001000100000:	sigmoid_prime = 18'b001100001101110011;
		14'b00001000100001:	sigmoid_prime = 18'b001100001101000011;
		14'b00001000100010:	sigmoid_prime = 18'b001100001100010100;
		14'b00001000100011:	sigmoid_prime = 18'b001100001011100100;
		14'b00001000100100:	sigmoid_prime = 18'b001100001010110100;
		14'b00001000100101:	sigmoid_prime = 18'b001100001010000101;
		14'b00001000100110:	sigmoid_prime = 18'b001100001001010101;
		14'b00001000100111:	sigmoid_prime = 18'b001100001000100101;
		14'b00001000101000:	sigmoid_prime = 18'b001100000111110110;
		14'b00001000101001:	sigmoid_prime = 18'b001100000111000110;
		14'b00001000101010:	sigmoid_prime = 18'b001100000110010110;
		14'b00001000101011:	sigmoid_prime = 18'b001100000101100110;
		14'b00001000101100:	sigmoid_prime = 18'b001100000100110110;
		14'b00001000101101:	sigmoid_prime = 18'b001100000100000111;
		14'b00001000101110:	sigmoid_prime = 18'b001100000011010111;
		14'b00001000101111:	sigmoid_prime = 18'b001100000010100111;
		14'b00001000110000:	sigmoid_prime = 18'b001100000001110111;
		14'b00001000110001:	sigmoid_prime = 18'b001100000001000111;
		14'b00001000110010:	sigmoid_prime = 18'b001100000000010111;
		14'b00001000110011:	sigmoid_prime = 18'b001011111111100111;
		14'b00001000110100:	sigmoid_prime = 18'b001011111110110111;
		14'b00001000110101:	sigmoid_prime = 18'b001011111110000111;
		14'b00001000110110:	sigmoid_prime = 18'b001011111101010111;
		14'b00001000110111:	sigmoid_prime = 18'b001011111100100111;
		14'b00001000111000:	sigmoid_prime = 18'b001011111011110111;
		14'b00001000111001:	sigmoid_prime = 18'b001011111011000111;
		14'b00001000111010:	sigmoid_prime = 18'b001011111010010110;
		14'b00001000111011:	sigmoid_prime = 18'b001011111001100110;
		14'b00001000111100:	sigmoid_prime = 18'b001011111000110110;
		14'b00001000111101:	sigmoid_prime = 18'b001011111000000110;
		14'b00001000111110:	sigmoid_prime = 18'b001011110111010110;
		14'b00001000111111:	sigmoid_prime = 18'b001011110110100101;
		14'b00001001000000:	sigmoid_prime = 18'b001011110101110101;
		14'b00001001000001:	sigmoid_prime = 18'b001011110101000101;
		14'b00001001000010:	sigmoid_prime = 18'b001011110100010100;
		14'b00001001000011:	sigmoid_prime = 18'b001011110011100100;
		14'b00001001000100:	sigmoid_prime = 18'b001011110010110100;
		14'b00001001000101:	sigmoid_prime = 18'b001011110010000011;
		14'b00001001000110:	sigmoid_prime = 18'b001011110001010011;
		14'b00001001000111:	sigmoid_prime = 18'b001011110000100010;
		14'b00001001001000:	sigmoid_prime = 18'b001011101111110010;
		14'b00001001001001:	sigmoid_prime = 18'b001011101111000001;
		14'b00001001001010:	sigmoid_prime = 18'b001011101110010001;
		14'b00001001001011:	sigmoid_prime = 18'b001011101101100001;
		14'b00001001001100:	sigmoid_prime = 18'b001011101100110000;
		14'b00001001001101:	sigmoid_prime = 18'b001011101011111111;
		14'b00001001001110:	sigmoid_prime = 18'b001011101011001111;
		14'b00001001001111:	sigmoid_prime = 18'b001011101010011110;
		14'b00001001010000:	sigmoid_prime = 18'b001011101001101110;
		14'b00001001010001:	sigmoid_prime = 18'b001011101000111101;
		14'b00001001010010:	sigmoid_prime = 18'b001011101000001101;
		14'b00001001010011:	sigmoid_prime = 18'b001011100111011100;
		14'b00001001010100:	sigmoid_prime = 18'b001011100110101011;
		14'b00001001010101:	sigmoid_prime = 18'b001011100101111011;
		14'b00001001010110:	sigmoid_prime = 18'b001011100101001010;
		14'b00001001010111:	sigmoid_prime = 18'b001011100100011001;
		14'b00001001011000:	sigmoid_prime = 18'b001011100011101000;
		14'b00001001011001:	sigmoid_prime = 18'b001011100010111000;
		14'b00001001011010:	sigmoid_prime = 18'b001011100010000111;
		14'b00001001011011:	sigmoid_prime = 18'b001011100001010110;
		14'b00001001011100:	sigmoid_prime = 18'b001011100000100101;
		14'b00001001011101:	sigmoid_prime = 18'b001011011111110101;
		14'b00001001011110:	sigmoid_prime = 18'b001011011111000100;
		14'b00001001011111:	sigmoid_prime = 18'b001011011110010011;
		14'b00001001100000:	sigmoid_prime = 18'b001011011101100010;
		14'b00001001100001:	sigmoid_prime = 18'b001011011100110001;
		14'b00001001100010:	sigmoid_prime = 18'b001011011100000001;
		14'b00001001100011:	sigmoid_prime = 18'b001011011011010000;
		14'b00001001100100:	sigmoid_prime = 18'b001011011010011111;
		14'b00001001100101:	sigmoid_prime = 18'b001011011001101110;
		14'b00001001100110:	sigmoid_prime = 18'b001011011000111101;
		14'b00001001100111:	sigmoid_prime = 18'b001011011000001100;
		14'b00001001101000:	sigmoid_prime = 18'b001011010111011011;
		14'b00001001101001:	sigmoid_prime = 18'b001011010110101010;
		14'b00001001101010:	sigmoid_prime = 18'b001011010101111001;
		14'b00001001101011:	sigmoid_prime = 18'b001011010101001000;
		14'b00001001101100:	sigmoid_prime = 18'b001011010100010111;
		14'b00001001101101:	sigmoid_prime = 18'b001011010011100110;
		14'b00001001101110:	sigmoid_prime = 18'b001011010010110101;
		14'b00001001101111:	sigmoid_prime = 18'b001011010010000100;
		14'b00001001110000:	sigmoid_prime = 18'b001011010001010011;
		14'b00001001110001:	sigmoid_prime = 18'b001011010000100010;
		14'b00001001110010:	sigmoid_prime = 18'b001011001111110001;
		14'b00001001110011:	sigmoid_prime = 18'b001011001111000000;
		14'b00001001110100:	sigmoid_prime = 18'b001011001110001111;
		14'b00001001110101:	sigmoid_prime = 18'b001011001101011110;
		14'b00001001110110:	sigmoid_prime = 18'b001011001100101101;
		14'b00001001110111:	sigmoid_prime = 18'b001011001011111100;
		14'b00001001111000:	sigmoid_prime = 18'b001011001011001011;
		14'b00001001111001:	sigmoid_prime = 18'b001011001010011010;
		14'b00001001111010:	sigmoid_prime = 18'b001011001001101001;
		14'b00001001111011:	sigmoid_prime = 18'b001011001000111000;
		14'b00001001111100:	sigmoid_prime = 18'b001011001000000110;
		14'b00001001111101:	sigmoid_prime = 18'b001011000111010101;
		14'b00001001111110:	sigmoid_prime = 18'b001011000110100100;
		14'b00001001111111:	sigmoid_prime = 18'b001011000101110011;
		14'b00001010000000:	sigmoid_prime = 18'b001011000101000010;
		14'b00001010000001:	sigmoid_prime = 18'b001011000100010001;
		14'b00001010000010:	sigmoid_prime = 18'b001011000011100000;
		14'b00001010000011:	sigmoid_prime = 18'b001011000010101110;
		14'b00001010000100:	sigmoid_prime = 18'b001011000001111101;
		14'b00001010000101:	sigmoid_prime = 18'b001011000001001100;
		14'b00001010000110:	sigmoid_prime = 18'b001011000000011011;
		14'b00001010000111:	sigmoid_prime = 18'b001010111111101010;
		14'b00001010001000:	sigmoid_prime = 18'b001010111110111000;
		14'b00001010001001:	sigmoid_prime = 18'b001010111110000111;
		14'b00001010001010:	sigmoid_prime = 18'b001010111101010110;
		14'b00001010001011:	sigmoid_prime = 18'b001010111100100101;
		14'b00001010001100:	sigmoid_prime = 18'b001010111011110100;
		14'b00001010001101:	sigmoid_prime = 18'b001010111011000010;
		14'b00001010001110:	sigmoid_prime = 18'b001010111010010001;
		14'b00001010001111:	sigmoid_prime = 18'b001010111001100000;
		14'b00001010010000:	sigmoid_prime = 18'b001010111000101111;
		14'b00001010010001:	sigmoid_prime = 18'b001010110111111101;
		14'b00001010010010:	sigmoid_prime = 18'b001010110111001100;
		14'b00001010010011:	sigmoid_prime = 18'b001010110110011011;
		14'b00001010010100:	sigmoid_prime = 18'b001010110101101010;
		14'b00001010010101:	sigmoid_prime = 18'b001010110100111000;
		14'b00001010010110:	sigmoid_prime = 18'b001010110100000111;
		14'b00001010010111:	sigmoid_prime = 18'b001010110011010110;
		14'b00001010011000:	sigmoid_prime = 18'b001010110010100101;
		14'b00001010011001:	sigmoid_prime = 18'b001010110001110011;
		14'b00001010011010:	sigmoid_prime = 18'b001010110001000010;
		14'b00001010011011:	sigmoid_prime = 18'b001010110000010001;
		14'b00001010011100:	sigmoid_prime = 18'b001010101111100000;
		14'b00001010011101:	sigmoid_prime = 18'b001010101110101110;
		14'b00001010011110:	sigmoid_prime = 18'b001010101101111101;
		14'b00001010011111:	sigmoid_prime = 18'b001010101101001100;
		14'b00001010100000:	sigmoid_prime = 18'b001010101100011011;
		14'b00001010100001:	sigmoid_prime = 18'b001010101011101001;
		14'b00001010100010:	sigmoid_prime = 18'b001010101010111000;
		14'b00001010100011:	sigmoid_prime = 18'b001010101010000111;
		14'b00001010100100:	sigmoid_prime = 18'b001010101001010110;
		14'b00001010100101:	sigmoid_prime = 18'b001010101000100100;
		14'b00001010100110:	sigmoid_prime = 18'b001010100111110011;
		14'b00001010100111:	sigmoid_prime = 18'b001010100111000010;
		14'b00001010101000:	sigmoid_prime = 18'b001010100110010000;
		14'b00001010101001:	sigmoid_prime = 18'b001010100101011111;
		14'b00001010101010:	sigmoid_prime = 18'b001010100100101110;
		14'b00001010101011:	sigmoid_prime = 18'b001010100011111101;
		14'b00001010101100:	sigmoid_prime = 18'b001010100011001011;
		14'b00001010101101:	sigmoid_prime = 18'b001010100010011010;
		14'b00001010101110:	sigmoid_prime = 18'b001010100001101001;
		14'b00001010101111:	sigmoid_prime = 18'b001010100000111000;
		14'b00001010110000:	sigmoid_prime = 18'b001010100000000110;
		14'b00001010110001:	sigmoid_prime = 18'b001010011111010101;
		14'b00001010110010:	sigmoid_prime = 18'b001010011110100100;
		14'b00001010110011:	sigmoid_prime = 18'b001010011101110011;
		14'b00001010110100:	sigmoid_prime = 18'b001010011101000001;
		14'b00001010110101:	sigmoid_prime = 18'b001010011100010000;
		14'b00001010110110:	sigmoid_prime = 18'b001010011011011111;
		14'b00001010110111:	sigmoid_prime = 18'b001010011010101110;
		14'b00001010111000:	sigmoid_prime = 18'b001010011001111101;
		14'b00001010111001:	sigmoid_prime = 18'b001010011001001011;
		14'b00001010111010:	sigmoid_prime = 18'b001010011000011010;
		14'b00001010111011:	sigmoid_prime = 18'b001010010111101001;
		14'b00001010111100:	sigmoid_prime = 18'b001010010110111000;
		14'b00001010111101:	sigmoid_prime = 18'b001010010110000110;
		14'b00001010111110:	sigmoid_prime = 18'b001010010101010101;
		14'b00001010111111:	sigmoid_prime = 18'b001010010100100100;
		14'b00001011000000:	sigmoid_prime = 18'b001010010011110011;
		14'b00001011000001:	sigmoid_prime = 18'b001010010011000010;
		14'b00001011000010:	sigmoid_prime = 18'b001010010010010001;
		14'b00001011000011:	sigmoid_prime = 18'b001010010001011111;
		14'b00001011000100:	sigmoid_prime = 18'b001010010000101110;
		14'b00001011000101:	sigmoid_prime = 18'b001010001111111101;
		14'b00001011000110:	sigmoid_prime = 18'b001010001111001100;
		14'b00001011000111:	sigmoid_prime = 18'b001010001110011011;
		14'b00001011001000:	sigmoid_prime = 18'b001010001101101010;
		14'b00001011001001:	sigmoid_prime = 18'b001010001100111000;
		14'b00001011001010:	sigmoid_prime = 18'b001010001100000111;
		14'b00001011001011:	sigmoid_prime = 18'b001010001011010110;
		14'b00001011001100:	sigmoid_prime = 18'b001010001010100101;
		14'b00001011001101:	sigmoid_prime = 18'b001010001001110100;
		14'b00001011001110:	sigmoid_prime = 18'b001010001001000011;
		14'b00001011001111:	sigmoid_prime = 18'b001010001000010010;
		14'b00001011010000:	sigmoid_prime = 18'b001010000111100001;
		14'b00001011010001:	sigmoid_prime = 18'b001010000110110000;
		14'b00001011010010:	sigmoid_prime = 18'b001010000101111111;
		14'b00001011010011:	sigmoid_prime = 18'b001010000101001110;
		14'b00001011010100:	sigmoid_prime = 18'b001010000100011100;
		14'b00001011010101:	sigmoid_prime = 18'b001010000011101011;
		14'b00001011010110:	sigmoid_prime = 18'b001010000010111010;
		14'b00001011010111:	sigmoid_prime = 18'b001010000010001001;
		14'b00001011011000:	sigmoid_prime = 18'b001010000001011000;
		14'b00001011011001:	sigmoid_prime = 18'b001010000000100111;
		14'b00001011011010:	sigmoid_prime = 18'b001001111111110110;
		14'b00001011011011:	sigmoid_prime = 18'b001001111111000101;
		14'b00001011011100:	sigmoid_prime = 18'b001001111110010100;
		14'b00001011011101:	sigmoid_prime = 18'b001001111101100011;
		14'b00001011011110:	sigmoid_prime = 18'b001001111100110010;
		14'b00001011011111:	sigmoid_prime = 18'b001001111100000010;
		14'b00001011100000:	sigmoid_prime = 18'b001001111011010001;
		14'b00001011100001:	sigmoid_prime = 18'b001001111010100000;
		14'b00001011100010:	sigmoid_prime = 18'b001001111001101111;
		14'b00001011100011:	sigmoid_prime = 18'b001001111000111110;
		14'b00001011100100:	sigmoid_prime = 18'b001001111000001101;
		14'b00001011100101:	sigmoid_prime = 18'b001001110111011100;
		14'b00001011100110:	sigmoid_prime = 18'b001001110110101011;
		14'b00001011100111:	sigmoid_prime = 18'b001001110101111010;
		14'b00001011101000:	sigmoid_prime = 18'b001001110101001010;
		14'b00001011101001:	sigmoid_prime = 18'b001001110100011001;
		14'b00001011101010:	sigmoid_prime = 18'b001001110011101000;
		14'b00001011101011:	sigmoid_prime = 18'b001001110010110111;
		14'b00001011101100:	sigmoid_prime = 18'b001001110010000110;
		14'b00001011101101:	sigmoid_prime = 18'b001001110001010110;
		14'b00001011101110:	sigmoid_prime = 18'b001001110000100101;
		14'b00001011101111:	sigmoid_prime = 18'b001001101111110100;
		14'b00001011110000:	sigmoid_prime = 18'b001001101111000011;
		14'b00001011110001:	sigmoid_prime = 18'b001001101110010011;
		14'b00001011110010:	sigmoid_prime = 18'b001001101101100010;
		14'b00001011110011:	sigmoid_prime = 18'b001001101100110001;
		14'b00001011110100:	sigmoid_prime = 18'b001001101100000000;
		14'b00001011110101:	sigmoid_prime = 18'b001001101011010000;
		14'b00001011110110:	sigmoid_prime = 18'b001001101010011111;
		14'b00001011110111:	sigmoid_prime = 18'b001001101001101110;
		14'b00001011111000:	sigmoid_prime = 18'b001001101000111110;
		14'b00001011111001:	sigmoid_prime = 18'b001001101000001101;
		14'b00001011111010:	sigmoid_prime = 18'b001001100111011101;
		14'b00001011111011:	sigmoid_prime = 18'b001001100110101100;
		14'b00001011111100:	sigmoid_prime = 18'b001001100101111011;
		14'b00001011111101:	sigmoid_prime = 18'b001001100101001011;
		14'b00001011111110:	sigmoid_prime = 18'b001001100100011010;
		14'b00001011111111:	sigmoid_prime = 18'b001001100011101010;
		14'b00001100000000:	sigmoid_prime = 18'b001001100010111001;
		14'b00001100000001:	sigmoid_prime = 18'b001001100010001001;
		14'b00001100000010:	sigmoid_prime = 18'b001001100001011000;
		14'b00001100000011:	sigmoid_prime = 18'b001001100000101000;
		14'b00001100000100:	sigmoid_prime = 18'b001001011111110111;
		14'b00001100000101:	sigmoid_prime = 18'b001001011111000111;
		14'b00001100000110:	sigmoid_prime = 18'b001001011110010111;
		14'b00001100000111:	sigmoid_prime = 18'b001001011101100110;
		14'b00001100001000:	sigmoid_prime = 18'b001001011100110110;
		14'b00001100001001:	sigmoid_prime = 18'b001001011100000101;
		14'b00001100001010:	sigmoid_prime = 18'b001001011011010101;
		14'b00001100001011:	sigmoid_prime = 18'b001001011010100101;
		14'b00001100001100:	sigmoid_prime = 18'b001001011001110100;
		14'b00001100001101:	sigmoid_prime = 18'b001001011001000100;
		14'b00001100001110:	sigmoid_prime = 18'b001001011000010100;
		14'b00001100001111:	sigmoid_prime = 18'b001001010111100100;
		14'b00001100010000:	sigmoid_prime = 18'b001001010110110011;
		14'b00001100010001:	sigmoid_prime = 18'b001001010110000011;
		14'b00001100010010:	sigmoid_prime = 18'b001001010101010011;
		14'b00001100010011:	sigmoid_prime = 18'b001001010100100011;
		14'b00001100010100:	sigmoid_prime = 18'b001001010011110011;
		14'b00001100010101:	sigmoid_prime = 18'b001001010011000010;
		14'b00001100010110:	sigmoid_prime = 18'b001001010010010010;
		14'b00001100010111:	sigmoid_prime = 18'b001001010001100010;
		14'b00001100011000:	sigmoid_prime = 18'b001001010000110010;
		14'b00001100011001:	sigmoid_prime = 18'b001001010000000010;
		14'b00001100011010:	sigmoid_prime = 18'b001001001111010010;
		14'b00001100011011:	sigmoid_prime = 18'b001001001110100010;
		14'b00001100011100:	sigmoid_prime = 18'b001001001101110010;
		14'b00001100011101:	sigmoid_prime = 18'b001001001101000010;
		14'b00001100011110:	sigmoid_prime = 18'b001001001100010010;
		14'b00001100011111:	sigmoid_prime = 18'b001001001011100010;
		14'b00001100100000:	sigmoid_prime = 18'b001001001010110010;
		14'b00001100100001:	sigmoid_prime = 18'b001001001010000010;
		14'b00001100100010:	sigmoid_prime = 18'b001001001001010010;
		14'b00001100100011:	sigmoid_prime = 18'b001001001000100010;
		14'b00001100100100:	sigmoid_prime = 18'b001001000111110011;
		14'b00001100100101:	sigmoid_prime = 18'b001001000111000011;
		14'b00001100100110:	sigmoid_prime = 18'b001001000110010011;
		14'b00001100100111:	sigmoid_prime = 18'b001001000101100011;
		14'b00001100101000:	sigmoid_prime = 18'b001001000100110011;
		14'b00001100101001:	sigmoid_prime = 18'b001001000100000100;
		14'b00001100101010:	sigmoid_prime = 18'b001001000011010100;
		14'b00001100101011:	sigmoid_prime = 18'b001001000010100100;
		14'b00001100101100:	sigmoid_prime = 18'b001001000001110100;
		14'b00001100101101:	sigmoid_prime = 18'b001001000001000101;
		14'b00001100101110:	sigmoid_prime = 18'b001001000000010101;
		14'b00001100101111:	sigmoid_prime = 18'b001000111111100110;
		14'b00001100110000:	sigmoid_prime = 18'b001000111110110110;
		14'b00001100110001:	sigmoid_prime = 18'b001000111110000110;
		14'b00001100110010:	sigmoid_prime = 18'b001000111101010111;
		14'b00001100110011:	sigmoid_prime = 18'b001000111100100111;
		14'b00001100110100:	sigmoid_prime = 18'b001000111011111000;
		14'b00001100110101:	sigmoid_prime = 18'b001000111011001000;
		14'b00001100110110:	sigmoid_prime = 18'b001000111010011001;
		14'b00001100110111:	sigmoid_prime = 18'b001000111001101001;
		14'b00001100111000:	sigmoid_prime = 18'b001000111000111010;
		14'b00001100111001:	sigmoid_prime = 18'b001000111000001011;
		14'b00001100111010:	sigmoid_prime = 18'b001000110111011011;
		14'b00001100111011:	sigmoid_prime = 18'b001000110110101100;
		14'b00001100111100:	sigmoid_prime = 18'b001000110101111100;
		14'b00001100111101:	sigmoid_prime = 18'b001000110101001101;
		14'b00001100111110:	sigmoid_prime = 18'b001000110100011110;
		14'b00001100111111:	sigmoid_prime = 18'b001000110011101111;
		14'b00001101000000:	sigmoid_prime = 18'b001000110010111111;
		14'b00001101000001:	sigmoid_prime = 18'b001000110010010000;
		14'b00001101000010:	sigmoid_prime = 18'b001000110001100001;
		14'b00001101000011:	sigmoid_prime = 18'b001000110000110010;
		14'b00001101000100:	sigmoid_prime = 18'b001000110000000011;
		14'b00001101000101:	sigmoid_prime = 18'b001000101111010100;
		14'b00001101000110:	sigmoid_prime = 18'b001000101110100101;
		14'b00001101000111:	sigmoid_prime = 18'b001000101101110101;
		14'b00001101001000:	sigmoid_prime = 18'b001000101101000110;
		14'b00001101001001:	sigmoid_prime = 18'b001000101100010111;
		14'b00001101001010:	sigmoid_prime = 18'b001000101011101000;
		14'b00001101001011:	sigmoid_prime = 18'b001000101010111001;
		14'b00001101001100:	sigmoid_prime = 18'b001000101010001011;
		14'b00001101001101:	sigmoid_prime = 18'b001000101001011100;
		14'b00001101001110:	sigmoid_prime = 18'b001000101000101101;
		14'b00001101001111:	sigmoid_prime = 18'b001000100111111110;
		14'b00001101010000:	sigmoid_prime = 18'b001000100111001111;
		14'b00001101010001:	sigmoid_prime = 18'b001000100110100000;
		14'b00001101010010:	sigmoid_prime = 18'b001000100101110001;
		14'b00001101010011:	sigmoid_prime = 18'b001000100101000011;
		14'b00001101010100:	sigmoid_prime = 18'b001000100100010100;
		14'b00001101010101:	sigmoid_prime = 18'b001000100011100101;
		14'b00001101010110:	sigmoid_prime = 18'b001000100010110111;
		14'b00001101010111:	sigmoid_prime = 18'b001000100010001000;
		14'b00001101011000:	sigmoid_prime = 18'b001000100001011001;
		14'b00001101011001:	sigmoid_prime = 18'b001000100000101011;
		14'b00001101011010:	sigmoid_prime = 18'b001000011111111100;
		14'b00001101011011:	sigmoid_prime = 18'b001000011111001110;
		14'b00001101011100:	sigmoid_prime = 18'b001000011110011111;
		14'b00001101011101:	sigmoid_prime = 18'b001000011101110001;
		14'b00001101011110:	sigmoid_prime = 18'b001000011101000010;
		14'b00001101011111:	sigmoid_prime = 18'b001000011100010100;
		14'b00001101100000:	sigmoid_prime = 18'b001000011011100101;
		14'b00001101100001:	sigmoid_prime = 18'b001000011010110111;
		14'b00001101100010:	sigmoid_prime = 18'b001000011010001001;
		14'b00001101100011:	sigmoid_prime = 18'b001000011001011010;
		14'b00001101100100:	sigmoid_prime = 18'b001000011000101100;
		14'b00001101100101:	sigmoid_prime = 18'b001000010111111110;
		14'b00001101100110:	sigmoid_prime = 18'b001000010111001111;
		14'b00001101100111:	sigmoid_prime = 18'b001000010110100001;
		14'b00001101101000:	sigmoid_prime = 18'b001000010101110011;
		14'b00001101101001:	sigmoid_prime = 18'b001000010101000101;
		14'b00001101101010:	sigmoid_prime = 18'b001000010100010111;
		14'b00001101101011:	sigmoid_prime = 18'b001000010011101001;
		14'b00001101101100:	sigmoid_prime = 18'b001000010010111011;
		14'b00001101101101:	sigmoid_prime = 18'b001000010010001101;
		14'b00001101101110:	sigmoid_prime = 18'b001000010001011111;
		14'b00001101101111:	sigmoid_prime = 18'b001000010000110001;
		14'b00001101110000:	sigmoid_prime = 18'b001000010000000011;
		14'b00001101110001:	sigmoid_prime = 18'b001000001111010101;
		14'b00001101110010:	sigmoid_prime = 18'b001000001110100111;
		14'b00001101110011:	sigmoid_prime = 18'b001000001101111001;
		14'b00001101110100:	sigmoid_prime = 18'b001000001101001011;
		14'b00001101110101:	sigmoid_prime = 18'b001000001100011101;
		14'b00001101110110:	sigmoid_prime = 18'b001000001011110000;
		14'b00001101110111:	sigmoid_prime = 18'b001000001011000010;
		14'b00001101111000:	sigmoid_prime = 18'b001000001010010100;
		14'b00001101111001:	sigmoid_prime = 18'b001000001001100110;
		14'b00001101111010:	sigmoid_prime = 18'b001000001000111001;
		14'b00001101111011:	sigmoid_prime = 18'b001000001000001011;
		14'b00001101111100:	sigmoid_prime = 18'b001000000111011110;
		14'b00001101111101:	sigmoid_prime = 18'b001000000110110000;
		14'b00001101111110:	sigmoid_prime = 18'b001000000110000010;
		14'b00001101111111:	sigmoid_prime = 18'b001000000101010101;
		14'b00001110000000:	sigmoid_prime = 18'b001000000100101000;
		14'b00001110000001:	sigmoid_prime = 18'b001000000011111010;
		14'b00001110000010:	sigmoid_prime = 18'b001000000011001101;
		14'b00001110000011:	sigmoid_prime = 18'b001000000010011111;
		14'b00001110000100:	sigmoid_prime = 18'b001000000001110010;
		14'b00001110000101:	sigmoid_prime = 18'b001000000001000101;
		14'b00001110000110:	sigmoid_prime = 18'b001000000000010111;
		14'b00001110000111:	sigmoid_prime = 18'b000111111111101010;
		14'b00001110001000:	sigmoid_prime = 18'b000111111110111101;
		14'b00001110001001:	sigmoid_prime = 18'b000111111110010000;
		14'b00001110001010:	sigmoid_prime = 18'b000111111101100010;
		14'b00001110001011:	sigmoid_prime = 18'b000111111100110101;
		14'b00001110001100:	sigmoid_prime = 18'b000111111100001000;
		14'b00001110001101:	sigmoid_prime = 18'b000111111011011011;
		14'b00001110001110:	sigmoid_prime = 18'b000111111010101110;
		14'b00001110001111:	sigmoid_prime = 18'b000111111010000001;
		14'b00001110010000:	sigmoid_prime = 18'b000111111001010100;
		14'b00001110010001:	sigmoid_prime = 18'b000111111000100111;
		14'b00001110010010:	sigmoid_prime = 18'b000111110111111010;
		14'b00001110010011:	sigmoid_prime = 18'b000111110111001101;
		14'b00001110010100:	sigmoid_prime = 18'b000111110110100001;
		14'b00001110010101:	sigmoid_prime = 18'b000111110101110100;
		14'b00001110010110:	sigmoid_prime = 18'b000111110101000111;
		14'b00001110010111:	sigmoid_prime = 18'b000111110100011010;
		14'b00001110011000:	sigmoid_prime = 18'b000111110011101110;
		14'b00001110011001:	sigmoid_prime = 18'b000111110011000001;
		14'b00001110011010:	sigmoid_prime = 18'b000111110010010100;
		14'b00001110011011:	sigmoid_prime = 18'b000111110001101000;
		14'b00001110011100:	sigmoid_prime = 18'b000111110000111011;
		14'b00001110011101:	sigmoid_prime = 18'b000111110000001111;
		14'b00001110011110:	sigmoid_prime = 18'b000111101111100010;
		14'b00001110011111:	sigmoid_prime = 18'b000111101110110110;
		14'b00001110100000:	sigmoid_prime = 18'b000111101110001001;
		14'b00001110100001:	sigmoid_prime = 18'b000111101101011101;
		14'b00001110100010:	sigmoid_prime = 18'b000111101100110000;
		14'b00001110100011:	sigmoid_prime = 18'b000111101100000100;
		14'b00001110100100:	sigmoid_prime = 18'b000111101011011000;
		14'b00001110100101:	sigmoid_prime = 18'b000111101010101011;
		14'b00001110100110:	sigmoid_prime = 18'b000111101001111111;
		14'b00001110100111:	sigmoid_prime = 18'b000111101001010011;
		14'b00001110101000:	sigmoid_prime = 18'b000111101000100111;
		14'b00001110101001:	sigmoid_prime = 18'b000111100111111011;
		14'b00001110101010:	sigmoid_prime = 18'b000111100111001110;
		14'b00001110101011:	sigmoid_prime = 18'b000111100110100010;
		14'b00001110101100:	sigmoid_prime = 18'b000111100101110110;
		14'b00001110101101:	sigmoid_prime = 18'b000111100101001010;
		14'b00001110101110:	sigmoid_prime = 18'b000111100100011110;
		14'b00001110101111:	sigmoid_prime = 18'b000111100011110010;
		14'b00001110110000:	sigmoid_prime = 18'b000111100011000110;
		14'b00001110110001:	sigmoid_prime = 18'b000111100010011011;
		14'b00001110110010:	sigmoid_prime = 18'b000111100001101111;
		14'b00001110110011:	sigmoid_prime = 18'b000111100001000011;
		14'b00001110110100:	sigmoid_prime = 18'b000111100000010111;
		14'b00001110110101:	sigmoid_prime = 18'b000111011111101011;
		14'b00001110110110:	sigmoid_prime = 18'b000111011111000000;
		14'b00001110110111:	sigmoid_prime = 18'b000111011110010100;
		14'b00001110111000:	sigmoid_prime = 18'b000111011101101000;
		14'b00001110111001:	sigmoid_prime = 18'b000111011100111101;
		14'b00001110111010:	sigmoid_prime = 18'b000111011100010001;
		14'b00001110111011:	sigmoid_prime = 18'b000111011011100110;
		14'b00001110111100:	sigmoid_prime = 18'b000111011010111010;
		14'b00001110111101:	sigmoid_prime = 18'b000111011010001111;
		14'b00001110111110:	sigmoid_prime = 18'b000111011001100011;
		14'b00001110111111:	sigmoid_prime = 18'b000111011000111000;
		14'b00001111000000:	sigmoid_prime = 18'b000111011000001101;
		14'b00001111000001:	sigmoid_prime = 18'b000111010111100001;
		14'b00001111000010:	sigmoid_prime = 18'b000111010110110110;
		14'b00001111000011:	sigmoid_prime = 18'b000111010110001011;
		14'b00001111000100:	sigmoid_prime = 18'b000111010101100000;
		14'b00001111000101:	sigmoid_prime = 18'b000111010100110101;
		14'b00001111000110:	sigmoid_prime = 18'b000111010100001001;
		14'b00001111000111:	sigmoid_prime = 18'b000111010011011110;
		14'b00001111001000:	sigmoid_prime = 18'b000111010010110011;
		14'b00001111001001:	sigmoid_prime = 18'b000111010010001000;
		14'b00001111001010:	sigmoid_prime = 18'b000111010001011101;
		14'b00001111001011:	sigmoid_prime = 18'b000111010000110010;
		14'b00001111001100:	sigmoid_prime = 18'b000111010000000111;
		14'b00001111001101:	sigmoid_prime = 18'b000111001111011100;
		14'b00001111001110:	sigmoid_prime = 18'b000111001110110010;
		14'b00001111001111:	sigmoid_prime = 18'b000111001110000111;
		14'b00001111010000:	sigmoid_prime = 18'b000111001101011100;
		14'b00001111010001:	sigmoid_prime = 18'b000111001100110001;
		14'b00001111010010:	sigmoid_prime = 18'b000111001100000111;
		14'b00001111010011:	sigmoid_prime = 18'b000111001011011100;
		14'b00001111010100:	sigmoid_prime = 18'b000111001010110001;
		14'b00001111010101:	sigmoid_prime = 18'b000111001010000111;
		14'b00001111010110:	sigmoid_prime = 18'b000111001001011100;
		14'b00001111010111:	sigmoid_prime = 18'b000111001000110010;
		14'b00001111011000:	sigmoid_prime = 18'b000111001000000111;
		14'b00001111011001:	sigmoid_prime = 18'b000111000111011101;
		14'b00001111011010:	sigmoid_prime = 18'b000111000110110010;
		14'b00001111011011:	sigmoid_prime = 18'b000111000110001000;
		14'b00001111011100:	sigmoid_prime = 18'b000111000101011110;
		14'b00001111011101:	sigmoid_prime = 18'b000111000100110011;
		14'b00001111011110:	sigmoid_prime = 18'b000111000100001001;
		14'b00001111011111:	sigmoid_prime = 18'b000111000011011111;
		14'b00001111100000:	sigmoid_prime = 18'b000111000010110101;
		14'b00001111100001:	sigmoid_prime = 18'b000111000010001011;
		14'b00001111100010:	sigmoid_prime = 18'b000111000001100000;
		14'b00001111100011:	sigmoid_prime = 18'b000111000000110110;
		14'b00001111100100:	sigmoid_prime = 18'b000111000000001100;
		14'b00001111100101:	sigmoid_prime = 18'b000110111111100010;
		14'b00001111100110:	sigmoid_prime = 18'b000110111110111000;
		14'b00001111100111:	sigmoid_prime = 18'b000110111110001110;
		14'b00001111101000:	sigmoid_prime = 18'b000110111101100101;
		14'b00001111101001:	sigmoid_prime = 18'b000110111100111011;
		14'b00001111101010:	sigmoid_prime = 18'b000110111100010001;
		14'b00001111101011:	sigmoid_prime = 18'b000110111011100111;
		14'b00001111101100:	sigmoid_prime = 18'b000110111010111101;
		14'b00001111101101:	sigmoid_prime = 18'b000110111010010100;
		14'b00001111101110:	sigmoid_prime = 18'b000110111001101010;
		14'b00001111101111:	sigmoid_prime = 18'b000110111001000001;
		14'b00001111110000:	sigmoid_prime = 18'b000110111000010111;
		14'b00001111110001:	sigmoid_prime = 18'b000110110111101101;
		14'b00001111110010:	sigmoid_prime = 18'b000110110111000100;
		14'b00001111110011:	sigmoid_prime = 18'b000110110110011010;
		14'b00001111110100:	sigmoid_prime = 18'b000110110101110001;
		14'b00001111110101:	sigmoid_prime = 18'b000110110101001000;
		14'b00001111110110:	sigmoid_prime = 18'b000110110100011110;
		14'b00001111110111:	sigmoid_prime = 18'b000110110011110101;
		14'b00001111111000:	sigmoid_prime = 18'b000110110011001100;
		14'b00001111111001:	sigmoid_prime = 18'b000110110010100010;
		14'b00001111111010:	sigmoid_prime = 18'b000110110001111001;
		14'b00001111111011:	sigmoid_prime = 18'b000110110001010000;
		14'b00001111111100:	sigmoid_prime = 18'b000110110000100111;
		14'b00001111111101:	sigmoid_prime = 18'b000110101111111110;
		14'b00001111111110:	sigmoid_prime = 18'b000110101111010101;
		14'b00001111111111:	sigmoid_prime = 18'b000110101110101100;
		14'b00010000000000:	sigmoid_prime = 18'b000110101110000011;
		14'b00010000000001:	sigmoid_prime = 18'b000110101101011010;
		14'b00010000000010:	sigmoid_prime = 18'b000110101100110001;
		14'b00010000000011:	sigmoid_prime = 18'b000110101100001000;
		14'b00010000000100:	sigmoid_prime = 18'b000110101011011111;
		14'b00010000000101:	sigmoid_prime = 18'b000110101010110111;
		14'b00010000000110:	sigmoid_prime = 18'b000110101010001110;
		14'b00010000000111:	sigmoid_prime = 18'b000110101001100101;
		14'b00010000001000:	sigmoid_prime = 18'b000110101000111101;
		14'b00010000001001:	sigmoid_prime = 18'b000110101000010100;
		14'b00010000001010:	sigmoid_prime = 18'b000110100111101011;
		14'b00010000001011:	sigmoid_prime = 18'b000110100111000011;
		14'b00010000001100:	sigmoid_prime = 18'b000110100110011010;
		14'b00010000001101:	sigmoid_prime = 18'b000110100101110010;
		14'b00010000001110:	sigmoid_prime = 18'b000110100101001010;
		14'b00010000001111:	sigmoid_prime = 18'b000110100100100001;
		14'b00010000010000:	sigmoid_prime = 18'b000110100011111001;
		14'b00010000010001:	sigmoid_prime = 18'b000110100011010001;
		14'b00010000010010:	sigmoid_prime = 18'b000110100010101000;
		14'b00010000010011:	sigmoid_prime = 18'b000110100010000000;
		14'b00010000010100:	sigmoid_prime = 18'b000110100001011000;
		14'b00010000010101:	sigmoid_prime = 18'b000110100000110000;
		14'b00010000010110:	sigmoid_prime = 18'b000110100000001000;
		14'b00010000010111:	sigmoid_prime = 18'b000110011111100000;
		14'b00010000011000:	sigmoid_prime = 18'b000110011110111000;
		14'b00010000011001:	sigmoid_prime = 18'b000110011110010000;
		14'b00010000011010:	sigmoid_prime = 18'b000110011101101000;
		14'b00010000011011:	sigmoid_prime = 18'b000110011101000000;
		14'b00010000011100:	sigmoid_prime = 18'b000110011100011000;
		14'b00010000011101:	sigmoid_prime = 18'b000110011011110000;
		14'b00010000011110:	sigmoid_prime = 18'b000110011011001000;
		14'b00010000011111:	sigmoid_prime = 18'b000110011010100001;
		14'b00010000100000:	sigmoid_prime = 18'b000110011001111001;
		14'b00010000100001:	sigmoid_prime = 18'b000110011001010001;
		14'b00010000100010:	sigmoid_prime = 18'b000110011000101010;
		14'b00010000100011:	sigmoid_prime = 18'b000110011000000010;
		14'b00010000100100:	sigmoid_prime = 18'b000110010111011011;
		14'b00010000100101:	sigmoid_prime = 18'b000110010110110011;
		14'b00010000100110:	sigmoid_prime = 18'b000110010110001100;
		14'b00010000100111:	sigmoid_prime = 18'b000110010101100100;
		14'b00010000101000:	sigmoid_prime = 18'b000110010100111101;
		14'b00010000101001:	sigmoid_prime = 18'b000110010100010101;
		14'b00010000101010:	sigmoid_prime = 18'b000110010011101110;
		14'b00010000101011:	sigmoid_prime = 18'b000110010011000111;
		14'b00010000101100:	sigmoid_prime = 18'b000110010010100000;
		14'b00010000101101:	sigmoid_prime = 18'b000110010001111001;
		14'b00010000101110:	sigmoid_prime = 18'b000110010001010001;
		14'b00010000101111:	sigmoid_prime = 18'b000110010000101010;
		14'b00010000110000:	sigmoid_prime = 18'b000110010000000011;
		14'b00010000110001:	sigmoid_prime = 18'b000110001111011100;
		14'b00010000110010:	sigmoid_prime = 18'b000110001110110101;
		14'b00010000110011:	sigmoid_prime = 18'b000110001110001110;
		14'b00010000110100:	sigmoid_prime = 18'b000110001101100111;
		14'b00010000110101:	sigmoid_prime = 18'b000110001101000001;
		14'b00010000110110:	sigmoid_prime = 18'b000110001100011010;
		14'b00010000110111:	sigmoid_prime = 18'b000110001011110011;
		14'b00010000111000:	sigmoid_prime = 18'b000110001011001100;
		14'b00010000111001:	sigmoid_prime = 18'b000110001010100110;
		14'b00010000111010:	sigmoid_prime = 18'b000110001001111111;
		14'b00010000111011:	sigmoid_prime = 18'b000110001001011000;
		14'b00010000111100:	sigmoid_prime = 18'b000110001000110010;
		14'b00010000111101:	sigmoid_prime = 18'b000110001000001011;
		14'b00010000111110:	sigmoid_prime = 18'b000110000111100101;
		14'b00010000111111:	sigmoid_prime = 18'b000110000110111110;
		14'b00010001000000:	sigmoid_prime = 18'b000110000110011000;
		14'b00010001000001:	sigmoid_prime = 18'b000110000101110001;
		14'b00010001000010:	sigmoid_prime = 18'b000110000101001011;
		14'b00010001000011:	sigmoid_prime = 18'b000110000100100101;
		14'b00010001000100:	sigmoid_prime = 18'b000110000011111111;
		14'b00010001000101:	sigmoid_prime = 18'b000110000011011000;
		14'b00010001000110:	sigmoid_prime = 18'b000110000010110010;
		14'b00010001000111:	sigmoid_prime = 18'b000110000010001100;
		14'b00010001001000:	sigmoid_prime = 18'b000110000001100110;
		14'b00010001001001:	sigmoid_prime = 18'b000110000001000000;
		14'b00010001001010:	sigmoid_prime = 18'b000110000000011010;
		14'b00010001001011:	sigmoid_prime = 18'b000101111111110100;
		14'b00010001001100:	sigmoid_prime = 18'b000101111111001110;
		14'b00010001001101:	sigmoid_prime = 18'b000101111110101000;
		14'b00010001001110:	sigmoid_prime = 18'b000101111110000010;
		14'b00010001001111:	sigmoid_prime = 18'b000101111101011101;
		14'b00010001010000:	sigmoid_prime = 18'b000101111100110111;
		14'b00010001010001:	sigmoid_prime = 18'b000101111100010001;
		14'b00010001010010:	sigmoid_prime = 18'b000101111011101100;
		14'b00010001010011:	sigmoid_prime = 18'b000101111011000110;
		14'b00010001010100:	sigmoid_prime = 18'b000101111010100000;
		14'b00010001010101:	sigmoid_prime = 18'b000101111001111011;
		14'b00010001010110:	sigmoid_prime = 18'b000101111001010101;
		14'b00010001010111:	sigmoid_prime = 18'b000101111000110000;
		14'b00010001011000:	sigmoid_prime = 18'b000101111000001010;
		14'b00010001011001:	sigmoid_prime = 18'b000101110111100101;
		14'b00010001011010:	sigmoid_prime = 18'b000101110111000000;
		14'b00010001011011:	sigmoid_prime = 18'b000101110110011010;
		14'b00010001011100:	sigmoid_prime = 18'b000101110101110101;
		14'b00010001011101:	sigmoid_prime = 18'b000101110101010000;
		14'b00010001011110:	sigmoid_prime = 18'b000101110100101011;
		14'b00010001011111:	sigmoid_prime = 18'b000101110100000110;
		14'b00010001100000:	sigmoid_prime = 18'b000101110011100001;
		14'b00010001100001:	sigmoid_prime = 18'b000101110010111011;
		14'b00010001100010:	sigmoid_prime = 18'b000101110010010110;
		14'b00010001100011:	sigmoid_prime = 18'b000101110001110001;
		14'b00010001100100:	sigmoid_prime = 18'b000101110001001101;
		14'b00010001100101:	sigmoid_prime = 18'b000101110000101000;
		14'b00010001100110:	sigmoid_prime = 18'b000101110000000011;
		14'b00010001100111:	sigmoid_prime = 18'b000101101111011110;
		14'b00010001101000:	sigmoid_prime = 18'b000101101110111001;
		14'b00010001101001:	sigmoid_prime = 18'b000101101110010101;
		14'b00010001101010:	sigmoid_prime = 18'b000101101101110000;
		14'b00010001101011:	sigmoid_prime = 18'b000101101101001011;
		14'b00010001101100:	sigmoid_prime = 18'b000101101100100111;
		14'b00010001101101:	sigmoid_prime = 18'b000101101100000010;
		14'b00010001101110:	sigmoid_prime = 18'b000101101011011110;
		14'b00010001101111:	sigmoid_prime = 18'b000101101010111001;
		14'b00010001110000:	sigmoid_prime = 18'b000101101010010101;
		14'b00010001110001:	sigmoid_prime = 18'b000101101001110000;
		14'b00010001110010:	sigmoid_prime = 18'b000101101001001100;
		14'b00010001110011:	sigmoid_prime = 18'b000101101000101000;
		14'b00010001110100:	sigmoid_prime = 18'b000101101000000011;
		14'b00010001110101:	sigmoid_prime = 18'b000101100111011111;
		14'b00010001110110:	sigmoid_prime = 18'b000101100110111011;
		14'b00010001110111:	sigmoid_prime = 18'b000101100110010111;
		14'b00010001111000:	sigmoid_prime = 18'b000101100101110011;
		14'b00010001111001:	sigmoid_prime = 18'b000101100101001111;
		14'b00010001111010:	sigmoid_prime = 18'b000101100100101011;
		14'b00010001111011:	sigmoid_prime = 18'b000101100100000111;
		14'b00010001111100:	sigmoid_prime = 18'b000101100011100011;
		14'b00010001111101:	sigmoid_prime = 18'b000101100010111111;
		14'b00010001111110:	sigmoid_prime = 18'b000101100010011011;
		14'b00010001111111:	sigmoid_prime = 18'b000101100001110111;
		14'b00010010000000:	sigmoid_prime = 18'b000101100001010100;
		14'b00010010000001:	sigmoid_prime = 18'b000101100000110000;
		14'b00010010000010:	sigmoid_prime = 18'b000101100000001100;
		14'b00010010000011:	sigmoid_prime = 18'b000101011111101000;
		14'b00010010000100:	sigmoid_prime = 18'b000101011111000101;
		14'b00010010000101:	sigmoid_prime = 18'b000101011110100001;
		14'b00010010000110:	sigmoid_prime = 18'b000101011101111110;
		14'b00010010000111:	sigmoid_prime = 18'b000101011101011010;
		14'b00010010001000:	sigmoid_prime = 18'b000101011100110111;
		14'b00010010001001:	sigmoid_prime = 18'b000101011100010100;
		14'b00010010001010:	sigmoid_prime = 18'b000101011011110000;
		14'b00010010001011:	sigmoid_prime = 18'b000101011011001101;
		14'b00010010001100:	sigmoid_prime = 18'b000101011010101010;
		14'b00010010001101:	sigmoid_prime = 18'b000101011010000110;
		14'b00010010001110:	sigmoid_prime = 18'b000101011001100011;
		14'b00010010001111:	sigmoid_prime = 18'b000101011001000000;
		14'b00010010010000:	sigmoid_prime = 18'b000101011000011101;
		14'b00010010010001:	sigmoid_prime = 18'b000101010111111010;
		14'b00010010010010:	sigmoid_prime = 18'b000101010111010111;
		14'b00010010010011:	sigmoid_prime = 18'b000101010110110100;
		14'b00010010010100:	sigmoid_prime = 18'b000101010110010001;
		14'b00010010010101:	sigmoid_prime = 18'b000101010101101110;
		14'b00010010010110:	sigmoid_prime = 18'b000101010101001011;
		14'b00010010010111:	sigmoid_prime = 18'b000101010100101000;
		14'b00010010011000:	sigmoid_prime = 18'b000101010100000110;
		14'b00010010011001:	sigmoid_prime = 18'b000101010011100011;
		14'b00010010011010:	sigmoid_prime = 18'b000101010011000000;
		14'b00010010011011:	sigmoid_prime = 18'b000101010010011110;
		14'b00010010011100:	sigmoid_prime = 18'b000101010001111011;
		14'b00010010011101:	sigmoid_prime = 18'b000101010001011000;
		14'b00010010011110:	sigmoid_prime = 18'b000101010000110110;
		14'b00010010011111:	sigmoid_prime = 18'b000101010000010100;
		14'b00010010100000:	sigmoid_prime = 18'b000101001111110001;
		14'b00010010100001:	sigmoid_prime = 18'b000101001111001111;
		14'b00010010100010:	sigmoid_prime = 18'b000101001110101100;
		14'b00010010100011:	sigmoid_prime = 18'b000101001110001010;
		14'b00010010100100:	sigmoid_prime = 18'b000101001101101000;
		14'b00010010100101:	sigmoid_prime = 18'b000101001101000110;
		14'b00010010100110:	sigmoid_prime = 18'b000101001100100011;
		14'b00010010100111:	sigmoid_prime = 18'b000101001100000001;
		14'b00010010101000:	sigmoid_prime = 18'b000101001011011111;
		14'b00010010101001:	sigmoid_prime = 18'b000101001010111101;
		14'b00010010101010:	sigmoid_prime = 18'b000101001010011011;
		14'b00010010101011:	sigmoid_prime = 18'b000101001001111001;
		14'b00010010101100:	sigmoid_prime = 18'b000101001001010111;
		14'b00010010101101:	sigmoid_prime = 18'b000101001000110101;
		14'b00010010101110:	sigmoid_prime = 18'b000101001000010011;
		14'b00010010101111:	sigmoid_prime = 18'b000101000111110010;
		14'b00010010110000:	sigmoid_prime = 18'b000101000111010000;
		14'b00010010110001:	sigmoid_prime = 18'b000101000110101110;
		14'b00010010110010:	sigmoid_prime = 18'b000101000110001100;
		14'b00010010110011:	sigmoid_prime = 18'b000101000101101011;
		14'b00010010110100:	sigmoid_prime = 18'b000101000101001001;
		14'b00010010110101:	sigmoid_prime = 18'b000101000100101000;
		14'b00010010110110:	sigmoid_prime = 18'b000101000100000110;
		14'b00010010110111:	sigmoid_prime = 18'b000101000011100101;
		14'b00010010111000:	sigmoid_prime = 18'b000101000011000011;
		14'b00010010111001:	sigmoid_prime = 18'b000101000010100010;
		14'b00010010111010:	sigmoid_prime = 18'b000101000010000001;
		14'b00010010111011:	sigmoid_prime = 18'b000101000001011111;
		14'b00010010111100:	sigmoid_prime = 18'b000101000000111110;
		14'b00010010111101:	sigmoid_prime = 18'b000101000000011101;
		14'b00010010111110:	sigmoid_prime = 18'b000100111111111100;
		14'b00010010111111:	sigmoid_prime = 18'b000100111111011010;
		14'b00010011000000:	sigmoid_prime = 18'b000100111110111001;
		14'b00010011000001:	sigmoid_prime = 18'b000100111110011000;
		14'b00010011000010:	sigmoid_prime = 18'b000100111101110111;
		14'b00010011000011:	sigmoid_prime = 18'b000100111101010110;
		14'b00010011000100:	sigmoid_prime = 18'b000100111100110101;
		14'b00010011000101:	sigmoid_prime = 18'b000100111100010100;
		14'b00010011000110:	sigmoid_prime = 18'b000100111011110100;
		14'b00010011000111:	sigmoid_prime = 18'b000100111011010011;
		14'b00010011001000:	sigmoid_prime = 18'b000100111010110010;
		14'b00010011001001:	sigmoid_prime = 18'b000100111010010001;
		14'b00010011001010:	sigmoid_prime = 18'b000100111001110001;
		14'b00010011001011:	sigmoid_prime = 18'b000100111001010000;
		14'b00010011001100:	sigmoid_prime = 18'b000100111000101111;
		14'b00010011001101:	sigmoid_prime = 18'b000100111000001111;
		14'b00010011001110:	sigmoid_prime = 18'b000100110111101110;
		14'b00010011001111:	sigmoid_prime = 18'b000100110111001110;
		14'b00010011010000:	sigmoid_prime = 18'b000100110110101101;
		14'b00010011010001:	sigmoid_prime = 18'b000100110110001101;
		14'b00010011010010:	sigmoid_prime = 18'b000100110101101101;
		14'b00010011010011:	sigmoid_prime = 18'b000100110101001100;
		14'b00010011010100:	sigmoid_prime = 18'b000100110100101100;
		14'b00010011010101:	sigmoid_prime = 18'b000100110100001100;
		14'b00010011010110:	sigmoid_prime = 18'b000100110011101100;
		14'b00010011010111:	sigmoid_prime = 18'b000100110011001011;
		14'b00010011011000:	sigmoid_prime = 18'b000100110010101011;
		14'b00010011011001:	sigmoid_prime = 18'b000100110010001011;
		14'b00010011011010:	sigmoid_prime = 18'b000100110001101011;
		14'b00010011011011:	sigmoid_prime = 18'b000100110001001011;
		14'b00010011011100:	sigmoid_prime = 18'b000100110000101011;
		14'b00010011011101:	sigmoid_prime = 18'b000100110000001011;
		14'b00010011011110:	sigmoid_prime = 18'b000100101111101100;
		14'b00010011011111:	sigmoid_prime = 18'b000100101111001100;
		14'b00010011100000:	sigmoid_prime = 18'b000100101110101100;
		14'b00010011100001:	sigmoid_prime = 18'b000100101110001100;
		14'b00010011100010:	sigmoid_prime = 18'b000100101101101101;
		14'b00010011100011:	sigmoid_prime = 18'b000100101101001101;
		14'b00010011100100:	sigmoid_prime = 18'b000100101100101101;
		14'b00010011100101:	sigmoid_prime = 18'b000100101100001110;
		14'b00010011100110:	sigmoid_prime = 18'b000100101011101110;
		14'b00010011100111:	sigmoid_prime = 18'b000100101011001111;
		14'b00010011101000:	sigmoid_prime = 18'b000100101010101111;
		14'b00010011101001:	sigmoid_prime = 18'b000100101010010000;
		14'b00010011101010:	sigmoid_prime = 18'b000100101001110000;
		14'b00010011101011:	sigmoid_prime = 18'b000100101001010001;
		14'b00010011101100:	sigmoid_prime = 18'b000100101000110010;
		14'b00010011101101:	sigmoid_prime = 18'b000100101000010011;
		14'b00010011101110:	sigmoid_prime = 18'b000100100111110011;
		14'b00010011101111:	sigmoid_prime = 18'b000100100111010100;
		14'b00010011110000:	sigmoid_prime = 18'b000100100110110101;
		14'b00010011110001:	sigmoid_prime = 18'b000100100110010110;
		14'b00010011110010:	sigmoid_prime = 18'b000100100101110111;
		14'b00010011110011:	sigmoid_prime = 18'b000100100101011000;
		14'b00010011110100:	sigmoid_prime = 18'b000100100100111001;
		14'b00010011110101:	sigmoid_prime = 18'b000100100100011010;
		14'b00010011110110:	sigmoid_prime = 18'b000100100011111011;
		14'b00010011110111:	sigmoid_prime = 18'b000100100011011100;
		14'b00010011111000:	sigmoid_prime = 18'b000100100010111110;
		14'b00010011111001:	sigmoid_prime = 18'b000100100010011111;
		14'b00010011111010:	sigmoid_prime = 18'b000100100010000000;
		14'b00010011111011:	sigmoid_prime = 18'b000100100001100010;
		14'b00010011111100:	sigmoid_prime = 18'b000100100001000011;
		14'b00010011111101:	sigmoid_prime = 18'b000100100000100100;
		14'b00010011111110:	sigmoid_prime = 18'b000100100000000110;
		14'b00010011111111:	sigmoid_prime = 18'b000100011111100111;
		14'b00010100000000:	sigmoid_prime = 18'b000100011111001001;
		14'b00010100000001:	sigmoid_prime = 18'b000100011110101010;
		14'b00010100000010:	sigmoid_prime = 18'b000100011110001100;
		14'b00010100000011:	sigmoid_prime = 18'b000100011101101110;
		14'b00010100000100:	sigmoid_prime = 18'b000100011101001111;
		14'b00010100000101:	sigmoid_prime = 18'b000100011100110001;
		14'b00010100000110:	sigmoid_prime = 18'b000100011100010011;
		14'b00010100000111:	sigmoid_prime = 18'b000100011011110101;
		14'b00010100001000:	sigmoid_prime = 18'b000100011011010110;
		14'b00010100001001:	sigmoid_prime = 18'b000100011010111000;
		14'b00010100001010:	sigmoid_prime = 18'b000100011010011010;
		14'b00010100001011:	sigmoid_prime = 18'b000100011001111100;
		14'b00010100001100:	sigmoid_prime = 18'b000100011001011110;
		14'b00010100001101:	sigmoid_prime = 18'b000100011001000000;
		14'b00010100001110:	sigmoid_prime = 18'b000100011000100010;
		14'b00010100001111:	sigmoid_prime = 18'b000100011000000101;
		14'b00010100010000:	sigmoid_prime = 18'b000100010111100111;
		14'b00010100010001:	sigmoid_prime = 18'b000100010111001001;
		14'b00010100010010:	sigmoid_prime = 18'b000100010110101011;
		14'b00010100010011:	sigmoid_prime = 18'b000100010110001110;
		14'b00010100010100:	sigmoid_prime = 18'b000100010101110000;
		14'b00010100010101:	sigmoid_prime = 18'b000100010101010010;
		14'b00010100010110:	sigmoid_prime = 18'b000100010100110101;
		14'b00010100010111:	sigmoid_prime = 18'b000100010100010111;
		14'b00010100011000:	sigmoid_prime = 18'b000100010011111010;
		14'b00010100011001:	sigmoid_prime = 18'b000100010011011100;
		14'b00010100011010:	sigmoid_prime = 18'b000100010010111111;
		14'b00010100011011:	sigmoid_prime = 18'b000100010010100001;
		14'b00010100011100:	sigmoid_prime = 18'b000100010010000100;
		14'b00010100011101:	sigmoid_prime = 18'b000100010001100111;
		14'b00010100011110:	sigmoid_prime = 18'b000100010001001010;
		14'b00010100011111:	sigmoid_prime = 18'b000100010000101100;
		14'b00010100100000:	sigmoid_prime = 18'b000100010000001111;
		14'b00010100100001:	sigmoid_prime = 18'b000100001111110010;
		14'b00010100100010:	sigmoid_prime = 18'b000100001111010101;
		14'b00010100100011:	sigmoid_prime = 18'b000100001110111000;
		14'b00010100100100:	sigmoid_prime = 18'b000100001110011011;
		14'b00010100100101:	sigmoid_prime = 18'b000100001101111110;
		14'b00010100100110:	sigmoid_prime = 18'b000100001101100001;
		14'b00010100100111:	sigmoid_prime = 18'b000100001101000100;
		14'b00010100101000:	sigmoid_prime = 18'b000100001100100111;
		14'b00010100101001:	sigmoid_prime = 18'b000100001100001010;
		14'b00010100101010:	sigmoid_prime = 18'b000100001011101110;
		14'b00010100101011:	sigmoid_prime = 18'b000100001011010001;
		14'b00010100101100:	sigmoid_prime = 18'b000100001010110100;
		14'b00010100101101:	sigmoid_prime = 18'b000100001010010111;
		14'b00010100101110:	sigmoid_prime = 18'b000100001001111011;
		14'b00010100101111:	sigmoid_prime = 18'b000100001001011110;
		14'b00010100110000:	sigmoid_prime = 18'b000100001001000010;
		14'b00010100110001:	sigmoid_prime = 18'b000100001000100101;
		14'b00010100110010:	sigmoid_prime = 18'b000100001000001001;
		14'b00010100110011:	sigmoid_prime = 18'b000100000111101100;
		14'b00010100110100:	sigmoid_prime = 18'b000100000111010000;
		14'b00010100110101:	sigmoid_prime = 18'b000100000110110100;
		14'b00010100110110:	sigmoid_prime = 18'b000100000110010111;
		14'b00010100110111:	sigmoid_prime = 18'b000100000101111011;
		14'b00010100111000:	sigmoid_prime = 18'b000100000101011111;
		14'b00010100111001:	sigmoid_prime = 18'b000100000101000011;
		14'b00010100111010:	sigmoid_prime = 18'b000100000100100110;
		14'b00010100111011:	sigmoid_prime = 18'b000100000100001010;
		14'b00010100111100:	sigmoid_prime = 18'b000100000011101110;
		14'b00010100111101:	sigmoid_prime = 18'b000100000011010010;
		14'b00010100111110:	sigmoid_prime = 18'b000100000010110110;
		14'b00010100111111:	sigmoid_prime = 18'b000100000010011010;
		14'b00010101000000:	sigmoid_prime = 18'b000100000001111110;
		14'b00010101000001:	sigmoid_prime = 18'b000100000001100011;
		14'b00010101000010:	sigmoid_prime = 18'b000100000001000111;
		14'b00010101000011:	sigmoid_prime = 18'b000100000000101011;
		14'b00010101000100:	sigmoid_prime = 18'b000100000000001111;
		14'b00010101000101:	sigmoid_prime = 18'b000011111111110011;
		14'b00010101000110:	sigmoid_prime = 18'b000011111111011000;
		14'b00010101000111:	sigmoid_prime = 18'b000011111110111100;
		14'b00010101001000:	sigmoid_prime = 18'b000011111110100001;
		14'b00010101001001:	sigmoid_prime = 18'b000011111110000101;
		14'b00010101001010:	sigmoid_prime = 18'b000011111101101001;
		14'b00010101001011:	sigmoid_prime = 18'b000011111101001110;
		14'b00010101001100:	sigmoid_prime = 18'b000011111100110011;
		14'b00010101001101:	sigmoid_prime = 18'b000011111100010111;
		14'b00010101001110:	sigmoid_prime = 18'b000011111011111100;
		14'b00010101001111:	sigmoid_prime = 18'b000011111011100000;
		14'b00010101010000:	sigmoid_prime = 18'b000011111011000101;
		14'b00010101010001:	sigmoid_prime = 18'b000011111010101010;
		14'b00010101010010:	sigmoid_prime = 18'b000011111010001111;
		14'b00010101010011:	sigmoid_prime = 18'b000011111001110100;
		14'b00010101010100:	sigmoid_prime = 18'b000011111001011000;
		14'b00010101010101:	sigmoid_prime = 18'b000011111000111101;
		14'b00010101010110:	sigmoid_prime = 18'b000011111000100010;
		14'b00010101010111:	sigmoid_prime = 18'b000011111000000111;
		14'b00010101011000:	sigmoid_prime = 18'b000011110111101100;
		14'b00010101011001:	sigmoid_prime = 18'b000011110111010001;
		14'b00010101011010:	sigmoid_prime = 18'b000011110110110110;
		14'b00010101011011:	sigmoid_prime = 18'b000011110110011100;
		14'b00010101011100:	sigmoid_prime = 18'b000011110110000001;
		14'b00010101011101:	sigmoid_prime = 18'b000011110101100110;
		14'b00010101011110:	sigmoid_prime = 18'b000011110101001011;
		14'b00010101011111:	sigmoid_prime = 18'b000011110100110000;
		14'b00010101100000:	sigmoid_prime = 18'b000011110100010110;
		14'b00010101100001:	sigmoid_prime = 18'b000011110011111011;
		14'b00010101100010:	sigmoid_prime = 18'b000011110011100001;
		14'b00010101100011:	sigmoid_prime = 18'b000011110011000110;
		14'b00010101100100:	sigmoid_prime = 18'b000011110010101100;
		14'b00010101100101:	sigmoid_prime = 18'b000011110010010001;
		14'b00010101100110:	sigmoid_prime = 18'b000011110001110111;
		14'b00010101100111:	sigmoid_prime = 18'b000011110001011100;
		14'b00010101101000:	sigmoid_prime = 18'b000011110001000010;
		14'b00010101101001:	sigmoid_prime = 18'b000011110000100111;
		14'b00010101101010:	sigmoid_prime = 18'b000011110000001101;
		14'b00010101101011:	sigmoid_prime = 18'b000011101111110011;
		14'b00010101101100:	sigmoid_prime = 18'b000011101111011001;
		14'b00010101101101:	sigmoid_prime = 18'b000011101110111111;
		14'b00010101101110:	sigmoid_prime = 18'b000011101110100100;
		14'b00010101101111:	sigmoid_prime = 18'b000011101110001010;
		14'b00010101110000:	sigmoid_prime = 18'b000011101101110000;
		14'b00010101110001:	sigmoid_prime = 18'b000011101101010110;
		14'b00010101110010:	sigmoid_prime = 18'b000011101100111100;
		14'b00010101110011:	sigmoid_prime = 18'b000011101100100010;
		14'b00010101110100:	sigmoid_prime = 18'b000011101100001000;
		14'b00010101110101:	sigmoid_prime = 18'b000011101011101111;
		14'b00010101110110:	sigmoid_prime = 18'b000011101011010101;
		14'b00010101110111:	sigmoid_prime = 18'b000011101010111011;
		14'b00010101111000:	sigmoid_prime = 18'b000011101010100001;
		14'b00010101111001:	sigmoid_prime = 18'b000011101010000111;
		14'b00010101111010:	sigmoid_prime = 18'b000011101001101110;
		14'b00010101111011:	sigmoid_prime = 18'b000011101001010100;
		14'b00010101111100:	sigmoid_prime = 18'b000011101000111010;
		14'b00010101111101:	sigmoid_prime = 18'b000011101000100001;
		14'b00010101111110:	sigmoid_prime = 18'b000011101000000111;
		14'b00010101111111:	sigmoid_prime = 18'b000011100111101110;
		14'b00010110000000:	sigmoid_prime = 18'b000011100111010100;
		14'b00010110000001:	sigmoid_prime = 18'b000011100110111011;
		14'b00010110000010:	sigmoid_prime = 18'b000011100110100010;
		14'b00010110000011:	sigmoid_prime = 18'b000011100110001000;
		14'b00010110000100:	sigmoid_prime = 18'b000011100101101111;
		14'b00010110000101:	sigmoid_prime = 18'b000011100101010110;
		14'b00010110000110:	sigmoid_prime = 18'b000011100100111100;
		14'b00010110000111:	sigmoid_prime = 18'b000011100100100011;
		14'b00010110001000:	sigmoid_prime = 18'b000011100100001010;
		14'b00010110001001:	sigmoid_prime = 18'b000011100011110001;
		14'b00010110001010:	sigmoid_prime = 18'b000011100011011000;
		14'b00010110001011:	sigmoid_prime = 18'b000011100010111111;
		14'b00010110001100:	sigmoid_prime = 18'b000011100010100110;
		14'b00010110001101:	sigmoid_prime = 18'b000011100010001101;
		14'b00010110001110:	sigmoid_prime = 18'b000011100001110100;
		14'b00010110001111:	sigmoid_prime = 18'b000011100001011011;
		14'b00010110010000:	sigmoid_prime = 18'b000011100001000010;
		14'b00010110010001:	sigmoid_prime = 18'b000011100000101001;
		14'b00010110010010:	sigmoid_prime = 18'b000011100000010000;
		14'b00010110010011:	sigmoid_prime = 18'b000011011111111000;
		14'b00010110010100:	sigmoid_prime = 18'b000011011111011111;
		14'b00010110010101:	sigmoid_prime = 18'b000011011111000110;
		14'b00010110010110:	sigmoid_prime = 18'b000011011110101110;
		14'b00010110010111:	sigmoid_prime = 18'b000011011110010101;
		14'b00010110011000:	sigmoid_prime = 18'b000011011101111101;
		14'b00010110011001:	sigmoid_prime = 18'b000011011101100100;
		14'b00010110011010:	sigmoid_prime = 18'b000011011101001011;
		14'b00010110011011:	sigmoid_prime = 18'b000011011100110011;
		14'b00010110011100:	sigmoid_prime = 18'b000011011100011011;
		14'b00010110011101:	sigmoid_prime = 18'b000011011100000010;
		14'b00010110011110:	sigmoid_prime = 18'b000011011011101010;
		14'b00010110011111:	sigmoid_prime = 18'b000011011011010010;
		14'b00010110100000:	sigmoid_prime = 18'b000011011010111001;
		14'b00010110100001:	sigmoid_prime = 18'b000011011010100001;
		14'b00010110100010:	sigmoid_prime = 18'b000011011010001001;
		14'b00010110100011:	sigmoid_prime = 18'b000011011001110001;
		14'b00010110100100:	sigmoid_prime = 18'b000011011001011000;
		14'b00010110100101:	sigmoid_prime = 18'b000011011001000000;
		14'b00010110100110:	sigmoid_prime = 18'b000011011000101000;
		14'b00010110100111:	sigmoid_prime = 18'b000011011000010000;
		14'b00010110101000:	sigmoid_prime = 18'b000011010111111000;
		14'b00010110101001:	sigmoid_prime = 18'b000011010111100000;
		14'b00010110101010:	sigmoid_prime = 18'b000011010111001000;
		14'b00010110101011:	sigmoid_prime = 18'b000011010110110001;
		14'b00010110101100:	sigmoid_prime = 18'b000011010110011001;
		14'b00010110101101:	sigmoid_prime = 18'b000011010110000001;
		14'b00010110101110:	sigmoid_prime = 18'b000011010101101001;
		14'b00010110101111:	sigmoid_prime = 18'b000011010101010001;
		14'b00010110110000:	sigmoid_prime = 18'b000011010100111010;
		14'b00010110110001:	sigmoid_prime = 18'b000011010100100010;
		14'b00010110110010:	sigmoid_prime = 18'b000011010100001010;
		14'b00010110110011:	sigmoid_prime = 18'b000011010011110011;
		14'b00010110110100:	sigmoid_prime = 18'b000011010011011011;
		14'b00010110110101:	sigmoid_prime = 18'b000011010011000100;
		14'b00010110110110:	sigmoid_prime = 18'b000011010010101100;
		14'b00010110110111:	sigmoid_prime = 18'b000011010010010101;
		14'b00010110111000:	sigmoid_prime = 18'b000011010001111101;
		14'b00010110111001:	sigmoid_prime = 18'b000011010001100110;
		14'b00010110111010:	sigmoid_prime = 18'b000011010001001111;
		14'b00010110111011:	sigmoid_prime = 18'b000011010000110111;
		14'b00010110111100:	sigmoid_prime = 18'b000011010000100000;
		14'b00010110111101:	sigmoid_prime = 18'b000011010000001001;
		14'b00010110111110:	sigmoid_prime = 18'b000011001111110010;
		14'b00010110111111:	sigmoid_prime = 18'b000011001111011010;
		14'b00010111000000:	sigmoid_prime = 18'b000011001111000011;
		14'b00010111000001:	sigmoid_prime = 18'b000011001110101100;
		14'b00010111000010:	sigmoid_prime = 18'b000011001110010101;
		14'b00010111000011:	sigmoid_prime = 18'b000011001101111110;
		14'b00010111000100:	sigmoid_prime = 18'b000011001101100111;
		14'b00010111000101:	sigmoid_prime = 18'b000011001101010000;
		14'b00010111000110:	sigmoid_prime = 18'b000011001100111001;
		14'b00010111000111:	sigmoid_prime = 18'b000011001100100010;
		14'b00010111001000:	sigmoid_prime = 18'b000011001100001011;
		14'b00010111001001:	sigmoid_prime = 18'b000011001011110101;
		14'b00010111001010:	sigmoid_prime = 18'b000011001011011110;
		14'b00010111001011:	sigmoid_prime = 18'b000011001011000111;
		14'b00010111001100:	sigmoid_prime = 18'b000011001010110000;
		14'b00010111001101:	sigmoid_prime = 18'b000011001010011010;
		14'b00010111001110:	sigmoid_prime = 18'b000011001010000011;
		14'b00010111001111:	sigmoid_prime = 18'b000011001001101100;
		14'b00010111010000:	sigmoid_prime = 18'b000011001001010110;
		14'b00010111010001:	sigmoid_prime = 18'b000011001000111111;
		14'b00010111010010:	sigmoid_prime = 18'b000011001000101001;
		14'b00010111010011:	sigmoid_prime = 18'b000011001000010010;
		14'b00010111010100:	sigmoid_prime = 18'b000011000111111100;
		14'b00010111010101:	sigmoid_prime = 18'b000011000111100101;
		14'b00010111010110:	sigmoid_prime = 18'b000011000111001111;
		14'b00010111010111:	sigmoid_prime = 18'b000011000110111001;
		14'b00010111011000:	sigmoid_prime = 18'b000011000110100010;
		14'b00010111011001:	sigmoid_prime = 18'b000011000110001100;
		14'b00010111011010:	sigmoid_prime = 18'b000011000101110110;
		14'b00010111011011:	sigmoid_prime = 18'b000011000101100000;
		14'b00010111011100:	sigmoid_prime = 18'b000011000101001010;
		14'b00010111011101:	sigmoid_prime = 18'b000011000100110011;
		14'b00010111011110:	sigmoid_prime = 18'b000011000100011101;
		14'b00010111011111:	sigmoid_prime = 18'b000011000100000111;
		14'b00010111100000:	sigmoid_prime = 18'b000011000011110001;
		14'b00010111100001:	sigmoid_prime = 18'b000011000011011011;
		14'b00010111100010:	sigmoid_prime = 18'b000011000011000101;
		14'b00010111100011:	sigmoid_prime = 18'b000011000010101111;
		14'b00010111100100:	sigmoid_prime = 18'b000011000010011010;
		14'b00010111100101:	sigmoid_prime = 18'b000011000010000100;
		14'b00010111100110:	sigmoid_prime = 18'b000011000001101110;
		14'b00010111100111:	sigmoid_prime = 18'b000011000001011000;
		14'b00010111101000:	sigmoid_prime = 18'b000011000001000010;
		14'b00010111101001:	sigmoid_prime = 18'b000011000000101101;
		14'b00010111101010:	sigmoid_prime = 18'b000011000000010111;
		14'b00010111101011:	sigmoid_prime = 18'b000011000000000001;
		14'b00010111101100:	sigmoid_prime = 18'b000010111111101100;
		14'b00010111101101:	sigmoid_prime = 18'b000010111111010110;
		14'b00010111101110:	sigmoid_prime = 18'b000010111111000001;
		14'b00010111101111:	sigmoid_prime = 18'b000010111110101011;
		14'b00010111110000:	sigmoid_prime = 18'b000010111110010110;
		14'b00010111110001:	sigmoid_prime = 18'b000010111110000000;
		14'b00010111110010:	sigmoid_prime = 18'b000010111101101011;
		14'b00010111110011:	sigmoid_prime = 18'b000010111101010101;
		14'b00010111110100:	sigmoid_prime = 18'b000010111101000000;
		14'b00010111110101:	sigmoid_prime = 18'b000010111100101011;
		14'b00010111110110:	sigmoid_prime = 18'b000010111100010101;
		14'b00010111110111:	sigmoid_prime = 18'b000010111100000000;
		14'b00010111111000:	sigmoid_prime = 18'b000010111011101011;
		14'b00010111111001:	sigmoid_prime = 18'b000010111011010110;
		14'b00010111111010:	sigmoid_prime = 18'b000010111011000001;
		14'b00010111111011:	sigmoid_prime = 18'b000010111010101011;
		14'b00010111111100:	sigmoid_prime = 18'b000010111010010110;
		14'b00010111111101:	sigmoid_prime = 18'b000010111010000001;
		14'b00010111111110:	sigmoid_prime = 18'b000010111001101100;
		14'b00010111111111:	sigmoid_prime = 18'b000010111001010111;
		14'b00011000000000:	sigmoid_prime = 18'b000010111001000010;
		14'b00011000000001:	sigmoid_prime = 18'b000010111000101101;
		14'b00011000000010:	sigmoid_prime = 18'b000010111000011000;
		14'b00011000000011:	sigmoid_prime = 18'b000010111000000100;
		14'b00011000000100:	sigmoid_prime = 18'b000010110111101111;
		14'b00011000000101:	sigmoid_prime = 18'b000010110111011010;
		14'b00011000000110:	sigmoid_prime = 18'b000010110111000101;
		14'b00011000000111:	sigmoid_prime = 18'b000010110110110001;
		14'b00011000001000:	sigmoid_prime = 18'b000010110110011100;
		14'b00011000001001:	sigmoid_prime = 18'b000010110110000111;
		14'b00011000001010:	sigmoid_prime = 18'b000010110101110011;
		14'b00011000001011:	sigmoid_prime = 18'b000010110101011110;
		14'b00011000001100:	sigmoid_prime = 18'b000010110101001001;
		14'b00011000001101:	sigmoid_prime = 18'b000010110100110101;
		14'b00011000001110:	sigmoid_prime = 18'b000010110100100000;
		14'b00011000001111:	sigmoid_prime = 18'b000010110100001100;
		14'b00011000010000:	sigmoid_prime = 18'b000010110011110111;
		14'b00011000010001:	sigmoid_prime = 18'b000010110011100011;
		14'b00011000010010:	sigmoid_prime = 18'b000010110011001111;
		14'b00011000010011:	sigmoid_prime = 18'b000010110010111010;
		14'b00011000010100:	sigmoid_prime = 18'b000010110010100110;
		14'b00011000010101:	sigmoid_prime = 18'b000010110010010010;
		14'b00011000010110:	sigmoid_prime = 18'b000010110001111110;
		14'b00011000010111:	sigmoid_prime = 18'b000010110001101001;
		14'b00011000011000:	sigmoid_prime = 18'b000010110001010101;
		14'b00011000011001:	sigmoid_prime = 18'b000010110001000001;
		14'b00011000011010:	sigmoid_prime = 18'b000010110000101101;
		14'b00011000011011:	sigmoid_prime = 18'b000010110000011001;
		14'b00011000011100:	sigmoid_prime = 18'b000010110000000101;
		14'b00011000011101:	sigmoid_prime = 18'b000010101111110001;
		14'b00011000011110:	sigmoid_prime = 18'b000010101111011101;
		14'b00011000011111:	sigmoid_prime = 18'b000010101111001001;
		14'b00011000100000:	sigmoid_prime = 18'b000010101110110101;
		14'b00011000100001:	sigmoid_prime = 18'b000010101110100001;
		14'b00011000100010:	sigmoid_prime = 18'b000010101110001101;
		14'b00011000100011:	sigmoid_prime = 18'b000010101101111001;
		14'b00011000100100:	sigmoid_prime = 18'b000010101101100110;
		14'b00011000100101:	sigmoid_prime = 18'b000010101101010010;
		14'b00011000100110:	sigmoid_prime = 18'b000010101100111110;
		14'b00011000100111:	sigmoid_prime = 18'b000010101100101010;
		14'b00011000101000:	sigmoid_prime = 18'b000010101100010111;
		14'b00011000101001:	sigmoid_prime = 18'b000010101100000011;
		14'b00011000101010:	sigmoid_prime = 18'b000010101011110000;
		14'b00011000101011:	sigmoid_prime = 18'b000010101011011100;
		14'b00011000101100:	sigmoid_prime = 18'b000010101011001000;
		14'b00011000101101:	sigmoid_prime = 18'b000010101010110101;
		14'b00011000101110:	sigmoid_prime = 18'b000010101010100001;
		14'b00011000101111:	sigmoid_prime = 18'b000010101010001110;
		14'b00011000110000:	sigmoid_prime = 18'b000010101001111011;
		14'b00011000110001:	sigmoid_prime = 18'b000010101001100111;
		14'b00011000110010:	sigmoid_prime = 18'b000010101001010100;
		14'b00011000110011:	sigmoid_prime = 18'b000010101001000001;
		14'b00011000110100:	sigmoid_prime = 18'b000010101000101101;
		14'b00011000110101:	sigmoid_prime = 18'b000010101000011010;
		14'b00011000110110:	sigmoid_prime = 18'b000010101000000111;
		14'b00011000110111:	sigmoid_prime = 18'b000010100111110100;
		14'b00011000111000:	sigmoid_prime = 18'b000010100111100000;
		14'b00011000111001:	sigmoid_prime = 18'b000010100111001101;
		14'b00011000111010:	sigmoid_prime = 18'b000010100110111010;
		14'b00011000111011:	sigmoid_prime = 18'b000010100110100111;
		14'b00011000111100:	sigmoid_prime = 18'b000010100110010100;
		14'b00011000111101:	sigmoid_prime = 18'b000010100110000001;
		14'b00011000111110:	sigmoid_prime = 18'b000010100101101110;
		14'b00011000111111:	sigmoid_prime = 18'b000010100101011011;
		14'b00011001000000:	sigmoid_prime = 18'b000010100101001000;
		14'b00011001000001:	sigmoid_prime = 18'b000010100100110101;
		14'b00011001000010:	sigmoid_prime = 18'b000010100100100010;
		14'b00011001000011:	sigmoid_prime = 18'b000010100100010000;
		14'b00011001000100:	sigmoid_prime = 18'b000010100011111101;
		14'b00011001000101:	sigmoid_prime = 18'b000010100011101010;
		14'b00011001000110:	sigmoid_prime = 18'b000010100011010111;
		14'b00011001000111:	sigmoid_prime = 18'b000010100011000101;
		14'b00011001001000:	sigmoid_prime = 18'b000010100010110010;
		14'b00011001001001:	sigmoid_prime = 18'b000010100010011111;
		14'b00011001001010:	sigmoid_prime = 18'b000010100010001101;
		14'b00011001001011:	sigmoid_prime = 18'b000010100001111010;
		14'b00011001001100:	sigmoid_prime = 18'b000010100001101000;
		14'b00011001001101:	sigmoid_prime = 18'b000010100001010101;
		14'b00011001001110:	sigmoid_prime = 18'b000010100001000011;
		14'b00011001001111:	sigmoid_prime = 18'b000010100000110000;
		14'b00011001010000:	sigmoid_prime = 18'b000010100000011110;
		14'b00011001010001:	sigmoid_prime = 18'b000010100000001011;
		14'b00011001010010:	sigmoid_prime = 18'b000010011111111001;
		14'b00011001010011:	sigmoid_prime = 18'b000010011111100110;
		14'b00011001010100:	sigmoid_prime = 18'b000010011111010100;
		14'b00011001010101:	sigmoid_prime = 18'b000010011111000010;
		14'b00011001010110:	sigmoid_prime = 18'b000010011110110000;
		14'b00011001010111:	sigmoid_prime = 18'b000010011110011101;
		14'b00011001011000:	sigmoid_prime = 18'b000010011110001011;
		14'b00011001011001:	sigmoid_prime = 18'b000010011101111001;
		14'b00011001011010:	sigmoid_prime = 18'b000010011101100111;
		14'b00011001011011:	sigmoid_prime = 18'b000010011101010101;
		14'b00011001011100:	sigmoid_prime = 18'b000010011101000011;
		14'b00011001011101:	sigmoid_prime = 18'b000010011100110001;
		14'b00011001011110:	sigmoid_prime = 18'b000010011100011111;
		14'b00011001011111:	sigmoid_prime = 18'b000010011100001101;
		14'b00011001100000:	sigmoid_prime = 18'b000010011011111011;
		14'b00011001100001:	sigmoid_prime = 18'b000010011011101001;
		14'b00011001100010:	sigmoid_prime = 18'b000010011011010111;
		14'b00011001100011:	sigmoid_prime = 18'b000010011011000101;
		14'b00011001100100:	sigmoid_prime = 18'b000010011010110011;
		14'b00011001100101:	sigmoid_prime = 18'b000010011010100001;
		14'b00011001100110:	sigmoid_prime = 18'b000010011010010000;
		14'b00011001100111:	sigmoid_prime = 18'b000010011001111110;
		14'b00011001101000:	sigmoid_prime = 18'b000010011001101100;
		14'b00011001101001:	sigmoid_prime = 18'b000010011001011010;
		14'b00011001101010:	sigmoid_prime = 18'b000010011001001001;
		14'b00011001101011:	sigmoid_prime = 18'b000010011000110111;
		14'b00011001101100:	sigmoid_prime = 18'b000010011000100101;
		14'b00011001101101:	sigmoid_prime = 18'b000010011000010100;
		14'b00011001101110:	sigmoid_prime = 18'b000010011000000010;
		14'b00011001101111:	sigmoid_prime = 18'b000010010111110001;
		14'b00011001110000:	sigmoid_prime = 18'b000010010111011111;
		14'b00011001110001:	sigmoid_prime = 18'b000010010111001110;
		14'b00011001110010:	sigmoid_prime = 18'b000010010110111100;
		14'b00011001110011:	sigmoid_prime = 18'b000010010110101011;
		14'b00011001110100:	sigmoid_prime = 18'b000010010110011010;
		14'b00011001110101:	sigmoid_prime = 18'b000010010110001000;
		14'b00011001110110:	sigmoid_prime = 18'b000010010101110111;
		14'b00011001110111:	sigmoid_prime = 18'b000010010101100110;
		14'b00011001111000:	sigmoid_prime = 18'b000010010101010100;
		14'b00011001111001:	sigmoid_prime = 18'b000010010101000011;
		14'b00011001111010:	sigmoid_prime = 18'b000010010100110010;
		14'b00011001111011:	sigmoid_prime = 18'b000010010100100001;
		14'b00011001111100:	sigmoid_prime = 18'b000010010100010000;
		14'b00011001111101:	sigmoid_prime = 18'b000010010011111110;
		14'b00011001111110:	sigmoid_prime = 18'b000010010011101101;
		14'b00011001111111:	sigmoid_prime = 18'b000010010011011100;
		14'b00011010000000:	sigmoid_prime = 18'b000010010011001011;
		14'b00011010000001:	sigmoid_prime = 18'b000010010010111010;
		14'b00011010000010:	sigmoid_prime = 18'b000010010010101001;
		14'b00011010000011:	sigmoid_prime = 18'b000010010010011000;
		14'b00011010000100:	sigmoid_prime = 18'b000010010010000111;
		14'b00011010000101:	sigmoid_prime = 18'b000010010001110111;
		14'b00011010000110:	sigmoid_prime = 18'b000010010001100110;
		14'b00011010000111:	sigmoid_prime = 18'b000010010001010101;
		14'b00011010001000:	sigmoid_prime = 18'b000010010001000100;
		14'b00011010001001:	sigmoid_prime = 18'b000010010000110011;
		14'b00011010001010:	sigmoid_prime = 18'b000010010000100010;
		14'b00011010001011:	sigmoid_prime = 18'b000010010000010010;
		14'b00011010001100:	sigmoid_prime = 18'b000010010000000001;
		14'b00011010001101:	sigmoid_prime = 18'b000010001111110000;
		14'b00011010001110:	sigmoid_prime = 18'b000010001111100000;
		14'b00011010001111:	sigmoid_prime = 18'b000010001111001111;
		14'b00011010010000:	sigmoid_prime = 18'b000010001110111110;
		14'b00011010010001:	sigmoid_prime = 18'b000010001110101110;
		14'b00011010010010:	sigmoid_prime = 18'b000010001110011101;
		14'b00011010010011:	sigmoid_prime = 18'b000010001110001101;
		14'b00011010010100:	sigmoid_prime = 18'b000010001101111100;
		14'b00011010010101:	sigmoid_prime = 18'b000010001101101100;
		14'b00011010010110:	sigmoid_prime = 18'b000010001101011011;
		14'b00011010010111:	sigmoid_prime = 18'b000010001101001011;
		14'b00011010011000:	sigmoid_prime = 18'b000010001100111011;
		14'b00011010011001:	sigmoid_prime = 18'b000010001100101010;
		14'b00011010011010:	sigmoid_prime = 18'b000010001100011010;
		14'b00011010011011:	sigmoid_prime = 18'b000010001100001010;
		14'b00011010011100:	sigmoid_prime = 18'b000010001011111010;
		14'b00011010011101:	sigmoid_prime = 18'b000010001011101001;
		14'b00011010011110:	sigmoid_prime = 18'b000010001011011001;
		14'b00011010011111:	sigmoid_prime = 18'b000010001011001001;
		14'b00011010100000:	sigmoid_prime = 18'b000010001010111001;
		14'b00011010100001:	sigmoid_prime = 18'b000010001010101001;
		14'b00011010100010:	sigmoid_prime = 18'b000010001010011000;
		14'b00011010100011:	sigmoid_prime = 18'b000010001010001000;
		14'b00011010100100:	sigmoid_prime = 18'b000010001001111000;
		14'b00011010100101:	sigmoid_prime = 18'b000010001001101000;
		14'b00011010100110:	sigmoid_prime = 18'b000010001001011000;
		14'b00011010100111:	sigmoid_prime = 18'b000010001001001000;
		14'b00011010101000:	sigmoid_prime = 18'b000010001000111000;
		14'b00011010101001:	sigmoid_prime = 18'b000010001000101001;
		14'b00011010101010:	sigmoid_prime = 18'b000010001000011001;
		14'b00011010101011:	sigmoid_prime = 18'b000010001000001001;
		14'b00011010101100:	sigmoid_prime = 18'b000010000111111001;
		14'b00011010101101:	sigmoid_prime = 18'b000010000111101001;
		14'b00011010101110:	sigmoid_prime = 18'b000010000111011001;
		14'b00011010101111:	sigmoid_prime = 18'b000010000111001010;
		14'b00011010110000:	sigmoid_prime = 18'b000010000110111010;
		14'b00011010110001:	sigmoid_prime = 18'b000010000110101010;
		14'b00011010110010:	sigmoid_prime = 18'b000010000110011011;
		14'b00011010110011:	sigmoid_prime = 18'b000010000110001011;
		14'b00011010110100:	sigmoid_prime = 18'b000010000101111011;
		14'b00011010110101:	sigmoid_prime = 18'b000010000101101100;
		14'b00011010110110:	sigmoid_prime = 18'b000010000101011100;
		14'b00011010110111:	sigmoid_prime = 18'b000010000101001101;
		14'b00011010111000:	sigmoid_prime = 18'b000010000100111101;
		14'b00011010111001:	sigmoid_prime = 18'b000010000100101110;
		14'b00011010111010:	sigmoid_prime = 18'b000010000100011110;
		14'b00011010111011:	sigmoid_prime = 18'b000010000100001111;
		14'b00011010111100:	sigmoid_prime = 18'b000010000011111111;
		14'b00011010111101:	sigmoid_prime = 18'b000010000011110000;
		14'b00011010111110:	sigmoid_prime = 18'b000010000011100000;
		14'b00011010111111:	sigmoid_prime = 18'b000010000011010001;
		14'b00011011000000:	sigmoid_prime = 18'b000010000011000010;
		14'b00011011000001:	sigmoid_prime = 18'b000010000010110011;
		14'b00011011000010:	sigmoid_prime = 18'b000010000010100011;
		14'b00011011000011:	sigmoid_prime = 18'b000010000010010100;
		14'b00011011000100:	sigmoid_prime = 18'b000010000010000101;
		14'b00011011000101:	sigmoid_prime = 18'b000010000001110110;
		14'b00011011000110:	sigmoid_prime = 18'b000010000001100111;
		14'b00011011000111:	sigmoid_prime = 18'b000010000001010111;
		14'b00011011001000:	sigmoid_prime = 18'b000010000001001000;
		14'b00011011001001:	sigmoid_prime = 18'b000010000000111001;
		14'b00011011001010:	sigmoid_prime = 18'b000010000000101010;
		14'b00011011001011:	sigmoid_prime = 18'b000010000000011011;
		14'b00011011001100:	sigmoid_prime = 18'b000010000000001100;
		14'b00011011001101:	sigmoid_prime = 18'b000001111111111101;
		14'b00011011001110:	sigmoid_prime = 18'b000001111111101110;
		14'b00011011001111:	sigmoid_prime = 18'b000001111111011111;
		14'b00011011010000:	sigmoid_prime = 18'b000001111111010000;
		14'b00011011010001:	sigmoid_prime = 18'b000001111111000010;
		14'b00011011010010:	sigmoid_prime = 18'b000001111110110011;
		14'b00011011010011:	sigmoid_prime = 18'b000001111110100100;
		14'b00011011010100:	sigmoid_prime = 18'b000001111110010101;
		14'b00011011010101:	sigmoid_prime = 18'b000001111110000110;
		14'b00011011010110:	sigmoid_prime = 18'b000001111101111000;
		14'b00011011010111:	sigmoid_prime = 18'b000001111101101001;
		14'b00011011011000:	sigmoid_prime = 18'b000001111101011010;
		14'b00011011011001:	sigmoid_prime = 18'b000001111101001011;
		14'b00011011011010:	sigmoid_prime = 18'b000001111100111101;
		14'b00011011011011:	sigmoid_prime = 18'b000001111100101110;
		14'b00011011011100:	sigmoid_prime = 18'b000001111100100000;
		14'b00011011011101:	sigmoid_prime = 18'b000001111100010001;
		14'b00011011011110:	sigmoid_prime = 18'b000001111100000010;
		14'b00011011011111:	sigmoid_prime = 18'b000001111011110100;
		14'b00011011100000:	sigmoid_prime = 18'b000001111011100101;
		14'b00011011100001:	sigmoid_prime = 18'b000001111011010111;
		14'b00011011100010:	sigmoid_prime = 18'b000001111011001000;
		14'b00011011100011:	sigmoid_prime = 18'b000001111010111010;
		14'b00011011100100:	sigmoid_prime = 18'b000001111010101100;
		14'b00011011100101:	sigmoid_prime = 18'b000001111010011101;
		14'b00011011100110:	sigmoid_prime = 18'b000001111010001111;
		14'b00011011100111:	sigmoid_prime = 18'b000001111010000001;
		14'b00011011101000:	sigmoid_prime = 18'b000001111001110010;
		14'b00011011101001:	sigmoid_prime = 18'b000001111001100100;
		14'b00011011101010:	sigmoid_prime = 18'b000001111001010110;
		14'b00011011101011:	sigmoid_prime = 18'b000001111001001000;
		14'b00011011101100:	sigmoid_prime = 18'b000001111000111001;
		14'b00011011101101:	sigmoid_prime = 18'b000001111000101011;
		14'b00011011101110:	sigmoid_prime = 18'b000001111000011101;
		14'b00011011101111:	sigmoid_prime = 18'b000001111000001111;
		14'b00011011110000:	sigmoid_prime = 18'b000001111000000001;
		14'b00011011110001:	sigmoid_prime = 18'b000001110111110011;
		14'b00011011110010:	sigmoid_prime = 18'b000001110111100101;
		14'b00011011110011:	sigmoid_prime = 18'b000001110111010111;
		14'b00011011110100:	sigmoid_prime = 18'b000001110111001001;
		14'b00011011110101:	sigmoid_prime = 18'b000001110110111011;
		14'b00011011110110:	sigmoid_prime = 18'b000001110110101101;
		14'b00011011110111:	sigmoid_prime = 18'b000001110110011111;
		14'b00011011111000:	sigmoid_prime = 18'b000001110110010001;
		14'b00011011111001:	sigmoid_prime = 18'b000001110110000011;
		14'b00011011111010:	sigmoid_prime = 18'b000001110101110101;
		14'b00011011111011:	sigmoid_prime = 18'b000001110101100111;
		14'b00011011111100:	sigmoid_prime = 18'b000001110101011001;
		14'b00011011111101:	sigmoid_prime = 18'b000001110101001100;
		14'b00011011111110:	sigmoid_prime = 18'b000001110100111110;
		14'b00011011111111:	sigmoid_prime = 18'b000001110100110000;
		14'b00011100000000:	sigmoid_prime = 18'b000001110100100010;
		14'b00011100000001:	sigmoid_prime = 18'b000001110100010101;
		14'b00011100000010:	sigmoid_prime = 18'b000001110100000111;
		14'b00011100000011:	sigmoid_prime = 18'b000001110011111001;
		14'b00011100000100:	sigmoid_prime = 18'b000001110011101100;
		14'b00011100000101:	sigmoid_prime = 18'b000001110011011110;
		14'b00011100000110:	sigmoid_prime = 18'b000001110011010000;
		14'b00011100000111:	sigmoid_prime = 18'b000001110011000011;
		14'b00011100001000:	sigmoid_prime = 18'b000001110010110101;
		14'b00011100001001:	sigmoid_prime = 18'b000001110010101000;
		14'b00011100001010:	sigmoid_prime = 18'b000001110010011010;
		14'b00011100001011:	sigmoid_prime = 18'b000001110010001101;
		14'b00011100001100:	sigmoid_prime = 18'b000001110001111111;
		14'b00011100001101:	sigmoid_prime = 18'b000001110001110010;
		14'b00011100001110:	sigmoid_prime = 18'b000001110001100101;
		14'b00011100001111:	sigmoid_prime = 18'b000001110001010111;
		14'b00011100010000:	sigmoid_prime = 18'b000001110001001010;
		14'b00011100010001:	sigmoid_prime = 18'b000001110000111101;
		14'b00011100010010:	sigmoid_prime = 18'b000001110000101111;
		14'b00011100010011:	sigmoid_prime = 18'b000001110000100010;
		14'b00011100010100:	sigmoid_prime = 18'b000001110000010101;
		14'b00011100010101:	sigmoid_prime = 18'b000001110000000111;
		14'b00011100010110:	sigmoid_prime = 18'b000001101111111010;
		14'b00011100010111:	sigmoid_prime = 18'b000001101111101101;
		14'b00011100011000:	sigmoid_prime = 18'b000001101111100000;
		14'b00011100011001:	sigmoid_prime = 18'b000001101111010011;
		14'b00011100011010:	sigmoid_prime = 18'b000001101111000110;
		14'b00011100011011:	sigmoid_prime = 18'b000001101110111001;
		14'b00011100011100:	sigmoid_prime = 18'b000001101110101011;
		14'b00011100011101:	sigmoid_prime = 18'b000001101110011110;
		14'b00011100011110:	sigmoid_prime = 18'b000001101110010001;
		14'b00011100011111:	sigmoid_prime = 18'b000001101110000100;
		14'b00011100100000:	sigmoid_prime = 18'b000001101101110111;
		14'b00011100100001:	sigmoid_prime = 18'b000001101101101010;
		14'b00011100100010:	sigmoid_prime = 18'b000001101101011101;
		14'b00011100100011:	sigmoid_prime = 18'b000001101101010001;
		14'b00011100100100:	sigmoid_prime = 18'b000001101101000100;
		14'b00011100100101:	sigmoid_prime = 18'b000001101100110111;
		14'b00011100100110:	sigmoid_prime = 18'b000001101100101010;
		14'b00011100100111:	sigmoid_prime = 18'b000001101100011101;
		14'b00011100101000:	sigmoid_prime = 18'b000001101100010000;
		14'b00011100101001:	sigmoid_prime = 18'b000001101100000011;
		14'b00011100101010:	sigmoid_prime = 18'b000001101011110111;
		14'b00011100101011:	sigmoid_prime = 18'b000001101011101010;
		14'b00011100101100:	sigmoid_prime = 18'b000001101011011101;
		14'b00011100101101:	sigmoid_prime = 18'b000001101011010001;
		14'b00011100101110:	sigmoid_prime = 18'b000001101011000100;
		14'b00011100101111:	sigmoid_prime = 18'b000001101010110111;
		14'b00011100110000:	sigmoid_prime = 18'b000001101010101011;
		14'b00011100110001:	sigmoid_prime = 18'b000001101010011110;
		14'b00011100110010:	sigmoid_prime = 18'b000001101010010001;
		14'b00011100110011:	sigmoid_prime = 18'b000001101010000101;
		14'b00011100110100:	sigmoid_prime = 18'b000001101001111000;
		14'b00011100110101:	sigmoid_prime = 18'b000001101001101100;
		14'b00011100110110:	sigmoid_prime = 18'b000001101001011111;
		14'b00011100110111:	sigmoid_prime = 18'b000001101001010011;
		14'b00011100111000:	sigmoid_prime = 18'b000001101001000110;
		14'b00011100111001:	sigmoid_prime = 18'b000001101000111010;
		14'b00011100111010:	sigmoid_prime = 18'b000001101000101101;
		14'b00011100111011:	sigmoid_prime = 18'b000001101000100001;
		14'b00011100111100:	sigmoid_prime = 18'b000001101000010101;
		14'b00011100111101:	sigmoid_prime = 18'b000001101000001000;
		14'b00011100111110:	sigmoid_prime = 18'b000001100111111100;
		14'b00011100111111:	sigmoid_prime = 18'b000001100111110000;
		14'b00011101000000:	sigmoid_prime = 18'b000001100111100011;
		14'b00011101000001:	sigmoid_prime = 18'b000001100111010111;
		14'b00011101000010:	sigmoid_prime = 18'b000001100111001011;
		14'b00011101000011:	sigmoid_prime = 18'b000001100110111111;
		14'b00011101000100:	sigmoid_prime = 18'b000001100110110011;
		14'b00011101000101:	sigmoid_prime = 18'b000001100110100110;
		14'b00011101000110:	sigmoid_prime = 18'b000001100110011010;
		14'b00011101000111:	sigmoid_prime = 18'b000001100110001110;
		14'b00011101001000:	sigmoid_prime = 18'b000001100110000010;
		14'b00011101001001:	sigmoid_prime = 18'b000001100101110110;
		14'b00011101001010:	sigmoid_prime = 18'b000001100101101010;
		14'b00011101001011:	sigmoid_prime = 18'b000001100101011110;
		14'b00011101001100:	sigmoid_prime = 18'b000001100101010010;
		14'b00011101001101:	sigmoid_prime = 18'b000001100101000110;
		14'b00011101001110:	sigmoid_prime = 18'b000001100100111010;
		14'b00011101001111:	sigmoid_prime = 18'b000001100100101110;
		14'b00011101010000:	sigmoid_prime = 18'b000001100100100010;
		14'b00011101010001:	sigmoid_prime = 18'b000001100100010110;
		14'b00011101010010:	sigmoid_prime = 18'b000001100100001010;
		14'b00011101010011:	sigmoid_prime = 18'b000001100011111110;
		14'b00011101010100:	sigmoid_prime = 18'b000001100011110010;
		14'b00011101010101:	sigmoid_prime = 18'b000001100011100110;
		14'b00011101010110:	sigmoid_prime = 18'b000001100011011011;
		14'b00011101010111:	sigmoid_prime = 18'b000001100011001111;
		14'b00011101011000:	sigmoid_prime = 18'b000001100011000011;
		14'b00011101011001:	sigmoid_prime = 18'b000001100010110111;
		14'b00011101011010:	sigmoid_prime = 18'b000001100010101011;
		14'b00011101011011:	sigmoid_prime = 18'b000001100010100000;
		14'b00011101011100:	sigmoid_prime = 18'b000001100010010100;
		14'b00011101011101:	sigmoid_prime = 18'b000001100010001000;
		14'b00011101011110:	sigmoid_prime = 18'b000001100001111101;
		14'b00011101011111:	sigmoid_prime = 18'b000001100001110001;
		14'b00011101100000:	sigmoid_prime = 18'b000001100001100110;
		14'b00011101100001:	sigmoid_prime = 18'b000001100001011010;
		14'b00011101100010:	sigmoid_prime = 18'b000001100001001110;
		14'b00011101100011:	sigmoid_prime = 18'b000001100001000011;
		14'b00011101100100:	sigmoid_prime = 18'b000001100000110111;
		14'b00011101100101:	sigmoid_prime = 18'b000001100000101100;
		14'b00011101100110:	sigmoid_prime = 18'b000001100000100000;
		14'b00011101100111:	sigmoid_prime = 18'b000001100000010101;
		14'b00011101101000:	sigmoid_prime = 18'b000001100000001001;
		14'b00011101101001:	sigmoid_prime = 18'b000001011111111110;
		14'b00011101101010:	sigmoid_prime = 18'b000001011111110010;
		14'b00011101101011:	sigmoid_prime = 18'b000001011111100111;
		14'b00011101101100:	sigmoid_prime = 18'b000001011111011100;
		14'b00011101101101:	sigmoid_prime = 18'b000001011111010000;
		14'b00011101101110:	sigmoid_prime = 18'b000001011111000101;
		14'b00011101101111:	sigmoid_prime = 18'b000001011110111010;
		14'b00011101110000:	sigmoid_prime = 18'b000001011110101110;
		14'b00011101110001:	sigmoid_prime = 18'b000001011110100011;
		14'b00011101110010:	sigmoid_prime = 18'b000001011110011000;
		14'b00011101110011:	sigmoid_prime = 18'b000001011110001101;
		14'b00011101110100:	sigmoid_prime = 18'b000001011110000001;
		14'b00011101110101:	sigmoid_prime = 18'b000001011101110110;
		14'b00011101110110:	sigmoid_prime = 18'b000001011101101011;
		14'b00011101110111:	sigmoid_prime = 18'b000001011101100000;
		14'b00011101111000:	sigmoid_prime = 18'b000001011101010101;
		14'b00011101111001:	sigmoid_prime = 18'b000001011101001010;
		14'b00011101111010:	sigmoid_prime = 18'b000001011100111111;
		14'b00011101111011:	sigmoid_prime = 18'b000001011100110100;
		14'b00011101111100:	sigmoid_prime = 18'b000001011100101000;
		14'b00011101111101:	sigmoid_prime = 18'b000001011100011101;
		14'b00011101111110:	sigmoid_prime = 18'b000001011100010010;
		14'b00011101111111:	sigmoid_prime = 18'b000001011100000111;
		14'b00011110000000:	sigmoid_prime = 18'b000001011011111100;
		14'b00011110000001:	sigmoid_prime = 18'b000001011011110010;
		14'b00011110000010:	sigmoid_prime = 18'b000001011011100111;
		14'b00011110000011:	sigmoid_prime = 18'b000001011011011100;
		14'b00011110000100:	sigmoid_prime = 18'b000001011011010001;
		14'b00011110000101:	sigmoid_prime = 18'b000001011011000110;
		14'b00011110000110:	sigmoid_prime = 18'b000001011010111011;
		14'b00011110000111:	sigmoid_prime = 18'b000001011010110000;
		14'b00011110001000:	sigmoid_prime = 18'b000001011010100101;
		14'b00011110001001:	sigmoid_prime = 18'b000001011010011011;
		14'b00011110001010:	sigmoid_prime = 18'b000001011010010000;
		14'b00011110001011:	sigmoid_prime = 18'b000001011010000101;
		14'b00011110001100:	sigmoid_prime = 18'b000001011001111010;
		14'b00011110001101:	sigmoid_prime = 18'b000001011001110000;
		14'b00011110001110:	sigmoid_prime = 18'b000001011001100101;
		14'b00011110001111:	sigmoid_prime = 18'b000001011001011010;
		14'b00011110010000:	sigmoid_prime = 18'b000001011001001111;
		14'b00011110010001:	sigmoid_prime = 18'b000001011001000101;
		14'b00011110010010:	sigmoid_prime = 18'b000001011000111010;
		14'b00011110010011:	sigmoid_prime = 18'b000001011000110000;
		14'b00011110010100:	sigmoid_prime = 18'b000001011000100101;
		14'b00011110010101:	sigmoid_prime = 18'b000001011000011010;
		14'b00011110010110:	sigmoid_prime = 18'b000001011000010000;
		14'b00011110010111:	sigmoid_prime = 18'b000001011000000101;
		14'b00011110011000:	sigmoid_prime = 18'b000001010111111011;
		14'b00011110011001:	sigmoid_prime = 18'b000001010111110000;
		14'b00011110011010:	sigmoid_prime = 18'b000001010111100110;
		14'b00011110011011:	sigmoid_prime = 18'b000001010111011011;
		14'b00011110011100:	sigmoid_prime = 18'b000001010111010001;
		14'b00011110011101:	sigmoid_prime = 18'b000001010111000111;
		14'b00011110011110:	sigmoid_prime = 18'b000001010110111100;
		14'b00011110011111:	sigmoid_prime = 18'b000001010110110010;
		14'b00011110100000:	sigmoid_prime = 18'b000001010110100111;
		14'b00011110100001:	sigmoid_prime = 18'b000001010110011101;
		14'b00011110100010:	sigmoid_prime = 18'b000001010110010011;
		14'b00011110100011:	sigmoid_prime = 18'b000001010110001000;
		14'b00011110100100:	sigmoid_prime = 18'b000001010101111110;
		14'b00011110100101:	sigmoid_prime = 18'b000001010101110100;
		14'b00011110100110:	sigmoid_prime = 18'b000001010101101010;
		14'b00011110100111:	sigmoid_prime = 18'b000001010101011111;
		14'b00011110101000:	sigmoid_prime = 18'b000001010101010101;
		14'b00011110101001:	sigmoid_prime = 18'b000001010101001011;
		14'b00011110101010:	sigmoid_prime = 18'b000001010101000001;
		14'b00011110101011:	sigmoid_prime = 18'b000001010100110111;
		14'b00011110101100:	sigmoid_prime = 18'b000001010100101100;
		14'b00011110101101:	sigmoid_prime = 18'b000001010100100010;
		14'b00011110101110:	sigmoid_prime = 18'b000001010100011000;
		14'b00011110101111:	sigmoid_prime = 18'b000001010100001110;
		14'b00011110110000:	sigmoid_prime = 18'b000001010100000100;
		14'b00011110110001:	sigmoid_prime = 18'b000001010011111010;
		14'b00011110110010:	sigmoid_prime = 18'b000001010011110000;
		14'b00011110110011:	sigmoid_prime = 18'b000001010011100110;
		14'b00011110110100:	sigmoid_prime = 18'b000001010011011100;
		14'b00011110110101:	sigmoid_prime = 18'b000001010011010010;
		14'b00011110110110:	sigmoid_prime = 18'b000001010011001000;
		14'b00011110110111:	sigmoid_prime = 18'b000001010010111110;
		14'b00011110111000:	sigmoid_prime = 18'b000001010010110100;
		14'b00011110111001:	sigmoid_prime = 18'b000001010010101010;
		14'b00011110111010:	sigmoid_prime = 18'b000001010010100000;
		14'b00011110111011:	sigmoid_prime = 18'b000001010010010110;
		14'b00011110111100:	sigmoid_prime = 18'b000001010010001100;
		14'b00011110111101:	sigmoid_prime = 18'b000001010010000011;
		14'b00011110111110:	sigmoid_prime = 18'b000001010001111001;
		14'b00011110111111:	sigmoid_prime = 18'b000001010001101111;
		14'b00011111000000:	sigmoid_prime = 18'b000001010001100101;
		14'b00011111000001:	sigmoid_prime = 18'b000001010001011011;
		14'b00011111000010:	sigmoid_prime = 18'b000001010001010010;
		14'b00011111000011:	sigmoid_prime = 18'b000001010001001000;
		14'b00011111000100:	sigmoid_prime = 18'b000001010000111110;
		14'b00011111000101:	sigmoid_prime = 18'b000001010000110100;
		14'b00011111000110:	sigmoid_prime = 18'b000001010000101011;
		14'b00011111000111:	sigmoid_prime = 18'b000001010000100001;
		14'b00011111001000:	sigmoid_prime = 18'b000001010000010111;
		14'b00011111001001:	sigmoid_prime = 18'b000001010000001110;
		14'b00011111001010:	sigmoid_prime = 18'b000001010000000100;
		14'b00011111001011:	sigmoid_prime = 18'b000001001111111011;
		14'b00011111001100:	sigmoid_prime = 18'b000001001111110001;
		14'b00011111001101:	sigmoid_prime = 18'b000001001111100111;
		14'b00011111001110:	sigmoid_prime = 18'b000001001111011110;
		14'b00011111001111:	sigmoid_prime = 18'b000001001111010100;
		14'b00011111010000:	sigmoid_prime = 18'b000001001111001011;
		14'b00011111010001:	sigmoid_prime = 18'b000001001111000001;
		14'b00011111010010:	sigmoid_prime = 18'b000001001110111000;
		14'b00011111010011:	sigmoid_prime = 18'b000001001110101110;
		14'b00011111010100:	sigmoid_prime = 18'b000001001110100101;
		14'b00011111010101:	sigmoid_prime = 18'b000001001110011011;
		14'b00011111010110:	sigmoid_prime = 18'b000001001110010010;
		14'b00011111010111:	sigmoid_prime = 18'b000001001110001001;
		14'b00011111011000:	sigmoid_prime = 18'b000001001101111111;
		14'b00011111011001:	sigmoid_prime = 18'b000001001101110110;
		14'b00011111011010:	sigmoid_prime = 18'b000001001101101101;
		14'b00011111011011:	sigmoid_prime = 18'b000001001101100011;
		14'b00011111011100:	sigmoid_prime = 18'b000001001101011010;
		14'b00011111011101:	sigmoid_prime = 18'b000001001101010001;
		14'b00011111011110:	sigmoid_prime = 18'b000001001101000111;
		14'b00011111011111:	sigmoid_prime = 18'b000001001100111110;
		14'b00011111100000:	sigmoid_prime = 18'b000001001100110101;
		14'b00011111100001:	sigmoid_prime = 18'b000001001100101100;
		14'b00011111100010:	sigmoid_prime = 18'b000001001100100010;
		14'b00011111100011:	sigmoid_prime = 18'b000001001100011001;
		14'b00011111100100:	sigmoid_prime = 18'b000001001100010000;
		14'b00011111100101:	sigmoid_prime = 18'b000001001100000111;
		14'b00011111100110:	sigmoid_prime = 18'b000001001011111110;
		14'b00011111100111:	sigmoid_prime = 18'b000001001011110101;
		14'b00011111101000:	sigmoid_prime = 18'b000001001011101100;
		14'b00011111101001:	sigmoid_prime = 18'b000001001011100010;
		14'b00011111101010:	sigmoid_prime = 18'b000001001011011001;
		14'b00011111101011:	sigmoid_prime = 18'b000001001011010000;
		14'b00011111101100:	sigmoid_prime = 18'b000001001011000111;
		14'b00011111101101:	sigmoid_prime = 18'b000001001010111110;
		14'b00011111101110:	sigmoid_prime = 18'b000001001010110101;
		14'b00011111101111:	sigmoid_prime = 18'b000001001010101100;
		14'b00011111110000:	sigmoid_prime = 18'b000001001010100011;
		14'b00011111110001:	sigmoid_prime = 18'b000001001010011010;
		14'b00011111110010:	sigmoid_prime = 18'b000001001010010001;
		14'b00011111110011:	sigmoid_prime = 18'b000001001010001000;
		14'b00011111110100:	sigmoid_prime = 18'b000001001001111111;
		14'b00011111110101:	sigmoid_prime = 18'b000001001001110111;
		14'b00011111110110:	sigmoid_prime = 18'b000001001001101110;
		14'b00011111110111:	sigmoid_prime = 18'b000001001001100101;
		14'b00011111111000:	sigmoid_prime = 18'b000001001001011100;
		14'b00011111111001:	sigmoid_prime = 18'b000001001001010011;
		14'b00011111111010:	sigmoid_prime = 18'b000001001001001010;
		14'b00011111111011:	sigmoid_prime = 18'b000001001001000001;
		14'b00011111111100:	sigmoid_prime = 18'b000001001000111001;
		14'b00011111111101:	sigmoid_prime = 18'b000001001000110000;
		14'b00011111111110:	sigmoid_prime = 18'b000001001000100111;
		14'b00011111111111:	sigmoid_prime = 18'b000001001000011110;
		14'b00100000000000:	sigmoid_prime = 18'b000001001000010110;
		14'b00100000000001:	sigmoid_prime = 18'b000001001000001101;
		14'b00100000000010:	sigmoid_prime = 18'b000001001000000100;
		14'b00100000000011:	sigmoid_prime = 18'b000001000111111100;
		14'b00100000000100:	sigmoid_prime = 18'b000001000111110011;
		14'b00100000000101:	sigmoid_prime = 18'b000001000111101010;
		14'b00100000000110:	sigmoid_prime = 18'b000001000111100010;
		14'b00100000000111:	sigmoid_prime = 18'b000001000111011001;
		14'b00100000001000:	sigmoid_prime = 18'b000001000111010000;
		14'b00100000001001:	sigmoid_prime = 18'b000001000111001000;
		14'b00100000001010:	sigmoid_prime = 18'b000001000110111111;
		14'b00100000001011:	sigmoid_prime = 18'b000001000110110111;
		14'b00100000001100:	sigmoid_prime = 18'b000001000110101110;
		14'b00100000001101:	sigmoid_prime = 18'b000001000110100110;
		14'b00100000001110:	sigmoid_prime = 18'b000001000110011101;
		14'b00100000001111:	sigmoid_prime = 18'b000001000110010101;
		14'b00100000010000:	sigmoid_prime = 18'b000001000110001100;
		14'b00100000010001:	sigmoid_prime = 18'b000001000110000100;
		14'b00100000010010:	sigmoid_prime = 18'b000001000101111011;
		14'b00100000010011:	sigmoid_prime = 18'b000001000101110011;
		14'b00100000010100:	sigmoid_prime = 18'b000001000101101010;
		14'b00100000010101:	sigmoid_prime = 18'b000001000101100010;
		14'b00100000010110:	sigmoid_prime = 18'b000001000101011010;
		14'b00100000010111:	sigmoid_prime = 18'b000001000101010001;
		14'b00100000011000:	sigmoid_prime = 18'b000001000101001001;
		14'b00100000011001:	sigmoid_prime = 18'b000001000101000001;
		14'b00100000011010:	sigmoid_prime = 18'b000001000100111000;
		14'b00100000011011:	sigmoid_prime = 18'b000001000100110000;
		14'b00100000011100:	sigmoid_prime = 18'b000001000100101000;
		14'b00100000011101:	sigmoid_prime = 18'b000001000100011111;
		14'b00100000011110:	sigmoid_prime = 18'b000001000100010111;
		14'b00100000011111:	sigmoid_prime = 18'b000001000100001111;
		14'b00100000100000:	sigmoid_prime = 18'b000001000100000111;
		14'b00100000100001:	sigmoid_prime = 18'b000001000011111110;
		14'b00100000100010:	sigmoid_prime = 18'b000001000011110110;
		14'b00100000100011:	sigmoid_prime = 18'b000001000011101110;
		14'b00100000100100:	sigmoid_prime = 18'b000001000011100110;
		14'b00100000100101:	sigmoid_prime = 18'b000001000011011110;
		14'b00100000100110:	sigmoid_prime = 18'b000001000011010110;
		14'b00100000100111:	sigmoid_prime = 18'b000001000011001101;
		14'b00100000101000:	sigmoid_prime = 18'b000001000011000101;
		14'b00100000101001:	sigmoid_prime = 18'b000001000010111101;
		14'b00100000101010:	sigmoid_prime = 18'b000001000010110101;
		14'b00100000101011:	sigmoid_prime = 18'b000001000010101101;
		14'b00100000101100:	sigmoid_prime = 18'b000001000010100101;
		14'b00100000101101:	sigmoid_prime = 18'b000001000010011101;
		14'b00100000101110:	sigmoid_prime = 18'b000001000010010101;
		14'b00100000101111:	sigmoid_prime = 18'b000001000010001101;
		14'b00100000110000:	sigmoid_prime = 18'b000001000010000101;
		14'b00100000110001:	sigmoid_prime = 18'b000001000001111101;
		14'b00100000110010:	sigmoid_prime = 18'b000001000001110101;
		14'b00100000110011:	sigmoid_prime = 18'b000001000001101101;
		14'b00100000110100:	sigmoid_prime = 18'b000001000001100101;
		14'b00100000110101:	sigmoid_prime = 18'b000001000001011101;
		14'b00100000110110:	sigmoid_prime = 18'b000001000001010101;
		14'b00100000110111:	sigmoid_prime = 18'b000001000001001101;
		14'b00100000111000:	sigmoid_prime = 18'b000001000001000101;
		14'b00100000111001:	sigmoid_prime = 18'b000001000000111110;
		14'b00100000111010:	sigmoid_prime = 18'b000001000000110110;
		14'b00100000111011:	sigmoid_prime = 18'b000001000000101110;
		14'b00100000111100:	sigmoid_prime = 18'b000001000000100110;
		14'b00100000111101:	sigmoid_prime = 18'b000001000000011110;
		14'b00100000111110:	sigmoid_prime = 18'b000001000000010110;
		14'b00100000111111:	sigmoid_prime = 18'b000001000000001111;
		14'b00100001000000:	sigmoid_prime = 18'b000001000000000111;
		14'b00100001000001:	sigmoid_prime = 18'b000000111111111111;
		14'b00100001000010:	sigmoid_prime = 18'b000000111111110111;
		14'b00100001000011:	sigmoid_prime = 18'b000000111111110000;
		14'b00100001000100:	sigmoid_prime = 18'b000000111111101000;
		14'b00100001000101:	sigmoid_prime = 18'b000000111111100000;
		14'b00100001000110:	sigmoid_prime = 18'b000000111111011001;
		14'b00100001000111:	sigmoid_prime = 18'b000000111111010001;
		14'b00100001001000:	sigmoid_prime = 18'b000000111111001001;
		14'b00100001001001:	sigmoid_prime = 18'b000000111111000010;
		14'b00100001001010:	sigmoid_prime = 18'b000000111110111010;
		14'b00100001001011:	sigmoid_prime = 18'b000000111110110010;
		14'b00100001001100:	sigmoid_prime = 18'b000000111110101011;
		14'b00100001001101:	sigmoid_prime = 18'b000000111110100011;
		14'b00100001001110:	sigmoid_prime = 18'b000000111110011100;
		14'b00100001001111:	sigmoid_prime = 18'b000000111110010100;
		14'b00100001010000:	sigmoid_prime = 18'b000000111110001101;
		14'b00100001010001:	sigmoid_prime = 18'b000000111110000101;
		14'b00100001010010:	sigmoid_prime = 18'b000000111101111110;
		14'b00100001010011:	sigmoid_prime = 18'b000000111101110110;
		14'b00100001010100:	sigmoid_prime = 18'b000000111101101111;
		14'b00100001010101:	sigmoid_prime = 18'b000000111101100111;
		14'b00100001010110:	sigmoid_prime = 18'b000000111101100000;
		14'b00100001010111:	sigmoid_prime = 18'b000000111101011000;
		14'b00100001011000:	sigmoid_prime = 18'b000000111101010001;
		14'b00100001011001:	sigmoid_prime = 18'b000000111101001001;
		14'b00100001011010:	sigmoid_prime = 18'b000000111101000010;
		14'b00100001011011:	sigmoid_prime = 18'b000000111100111011;
		14'b00100001011100:	sigmoid_prime = 18'b000000111100110011;
		14'b00100001011101:	sigmoid_prime = 18'b000000111100101100;
		14'b00100001011110:	sigmoid_prime = 18'b000000111100100100;
		14'b00100001011111:	sigmoid_prime = 18'b000000111100011101;
		14'b00100001100000:	sigmoid_prime = 18'b000000111100010110;
		14'b00100001100001:	sigmoid_prime = 18'b000000111100001110;
		14'b00100001100010:	sigmoid_prime = 18'b000000111100000111;
		14'b00100001100011:	sigmoid_prime = 18'b000000111100000000;
		14'b00100001100100:	sigmoid_prime = 18'b000000111011111001;
		14'b00100001100101:	sigmoid_prime = 18'b000000111011110001;
		14'b00100001100110:	sigmoid_prime = 18'b000000111011101010;
		14'b00100001100111:	sigmoid_prime = 18'b000000111011100011;
		14'b00100001101000:	sigmoid_prime = 18'b000000111011011100;
		14'b00100001101001:	sigmoid_prime = 18'b000000111011010100;
		14'b00100001101010:	sigmoid_prime = 18'b000000111011001101;
		14'b00100001101011:	sigmoid_prime = 18'b000000111011000110;
		14'b00100001101100:	sigmoid_prime = 18'b000000111010111111;
		14'b00100001101101:	sigmoid_prime = 18'b000000111010111000;
		14'b00100001101110:	sigmoid_prime = 18'b000000111010110001;
		14'b00100001101111:	sigmoid_prime = 18'b000000111010101001;
		14'b00100001110000:	sigmoid_prime = 18'b000000111010100010;
		14'b00100001110001:	sigmoid_prime = 18'b000000111010011011;
		14'b00100001110010:	sigmoid_prime = 18'b000000111010010100;
		14'b00100001110011:	sigmoid_prime = 18'b000000111010001101;
		14'b00100001110100:	sigmoid_prime = 18'b000000111010000110;
		14'b00100001110101:	sigmoid_prime = 18'b000000111001111111;
		14'b00100001110110:	sigmoid_prime = 18'b000000111001111000;
		14'b00100001110111:	sigmoid_prime = 18'b000000111001110001;
		14'b00100001111000:	sigmoid_prime = 18'b000000111001101010;
		14'b00100001111001:	sigmoid_prime = 18'b000000111001100011;
		14'b00100001111010:	sigmoid_prime = 18'b000000111001011100;
		14'b00100001111011:	sigmoid_prime = 18'b000000111001010101;
		14'b00100001111100:	sigmoid_prime = 18'b000000111001001110;
		14'b00100001111101:	sigmoid_prime = 18'b000000111001000111;
		14'b00100001111110:	sigmoid_prime = 18'b000000111001000000;
		14'b00100001111111:	sigmoid_prime = 18'b000000111000111001;
		14'b00100010000000:	sigmoid_prime = 18'b000000111000110010;
		14'b00100010000001:	sigmoid_prime = 18'b000000111000101011;
		14'b00100010000010:	sigmoid_prime = 18'b000000111000100101;
		14'b00100010000011:	sigmoid_prime = 18'b000000111000011110;
		14'b00100010000100:	sigmoid_prime = 18'b000000111000010111;
		14'b00100010000101:	sigmoid_prime = 18'b000000111000010000;
		14'b00100010000110:	sigmoid_prime = 18'b000000111000001001;
		14'b00100010000111:	sigmoid_prime = 18'b000000111000000010;
		14'b00100010001000:	sigmoid_prime = 18'b000000110111111100;
		14'b00100010001001:	sigmoid_prime = 18'b000000110111110101;
		14'b00100010001010:	sigmoid_prime = 18'b000000110111101110;
		14'b00100010001011:	sigmoid_prime = 18'b000000110111100111;
		14'b00100010001100:	sigmoid_prime = 18'b000000110111100000;
		14'b00100010001101:	sigmoid_prime = 18'b000000110111011010;
		14'b00100010001110:	sigmoid_prime = 18'b000000110111010011;
		14'b00100010001111:	sigmoid_prime = 18'b000000110111001100;
		14'b00100010010000:	sigmoid_prime = 18'b000000110111000110;
		14'b00100010010001:	sigmoid_prime = 18'b000000110110111111;
		14'b00100010010010:	sigmoid_prime = 18'b000000110110111000;
		14'b00100010010011:	sigmoid_prime = 18'b000000110110110010;
		14'b00100010010100:	sigmoid_prime = 18'b000000110110101011;
		14'b00100010010101:	sigmoid_prime = 18'b000000110110100100;
		14'b00100010010110:	sigmoid_prime = 18'b000000110110011110;
		14'b00100010010111:	sigmoid_prime = 18'b000000110110010111;
		14'b00100010011000:	sigmoid_prime = 18'b000000110110010000;
		14'b00100010011001:	sigmoid_prime = 18'b000000110110001010;
		14'b00100010011010:	sigmoid_prime = 18'b000000110110000011;
		14'b00100010011011:	sigmoid_prime = 18'b000000110101111101;
		14'b00100010011100:	sigmoid_prime = 18'b000000110101110110;
		14'b00100010011101:	sigmoid_prime = 18'b000000110101110000;
		14'b00100010011110:	sigmoid_prime = 18'b000000110101101001;
		14'b00100010011111:	sigmoid_prime = 18'b000000110101100010;
		14'b00100010100000:	sigmoid_prime = 18'b000000110101011100;
		14'b00100010100001:	sigmoid_prime = 18'b000000110101010101;
		14'b00100010100010:	sigmoid_prime = 18'b000000110101001111;
		14'b00100010100011:	sigmoid_prime = 18'b000000110101001000;
		14'b00100010100100:	sigmoid_prime = 18'b000000110101000010;
		14'b00100010100101:	sigmoid_prime = 18'b000000110100111100;
		14'b00100010100110:	sigmoid_prime = 18'b000000110100110101;
		14'b00100010100111:	sigmoid_prime = 18'b000000110100101111;
		14'b00100010101000:	sigmoid_prime = 18'b000000110100101000;
		14'b00100010101001:	sigmoid_prime = 18'b000000110100100010;
		14'b00100010101010:	sigmoid_prime = 18'b000000110100011100;
		14'b00100010101011:	sigmoid_prime = 18'b000000110100010101;
		14'b00100010101100:	sigmoid_prime = 18'b000000110100001111;
		14'b00100010101101:	sigmoid_prime = 18'b000000110100001000;
		14'b00100010101110:	sigmoid_prime = 18'b000000110100000010;
		14'b00100010101111:	sigmoid_prime = 18'b000000110011111100;
		14'b00100010110000:	sigmoid_prime = 18'b000000110011110101;
		14'b00100010110001:	sigmoid_prime = 18'b000000110011101111;
		14'b00100010110010:	sigmoid_prime = 18'b000000110011101001;
		14'b00100010110011:	sigmoid_prime = 18'b000000110011100011;
		14'b00100010110100:	sigmoid_prime = 18'b000000110011011100;
		14'b00100010110101:	sigmoid_prime = 18'b000000110011010110;
		14'b00100010110110:	sigmoid_prime = 18'b000000110011010000;
		14'b00100010110111:	sigmoid_prime = 18'b000000110011001001;
		14'b00100010111000:	sigmoid_prime = 18'b000000110011000011;
		14'b00100010111001:	sigmoid_prime = 18'b000000110010111101;
		14'b00100010111010:	sigmoid_prime = 18'b000000110010110111;
		14'b00100010111011:	sigmoid_prime = 18'b000000110010110001;
		14'b00100010111100:	sigmoid_prime = 18'b000000110010101010;
		14'b00100010111101:	sigmoid_prime = 18'b000000110010100100;
		14'b00100010111110:	sigmoid_prime = 18'b000000110010011110;
		14'b00100010111111:	sigmoid_prime = 18'b000000110010011000;
		14'b00100011000000:	sigmoid_prime = 18'b000000110010010010;
		14'b00100011000001:	sigmoid_prime = 18'b000000110010001100;
		14'b00100011000010:	sigmoid_prime = 18'b000000110010000110;
		14'b00100011000011:	sigmoid_prime = 18'b000000110010000000;
		14'b00100011000100:	sigmoid_prime = 18'b000000110001111001;
		14'b00100011000101:	sigmoid_prime = 18'b000000110001110011;
		14'b00100011000110:	sigmoid_prime = 18'b000000110001101101;
		14'b00100011000111:	sigmoid_prime = 18'b000000110001100111;
		14'b00100011001000:	sigmoid_prime = 18'b000000110001100001;
		14'b00100011001001:	sigmoid_prime = 18'b000000110001011011;
		14'b00100011001010:	sigmoid_prime = 18'b000000110001010101;
		14'b00100011001011:	sigmoid_prime = 18'b000000110001001111;
		14'b00100011001100:	sigmoid_prime = 18'b000000110001001001;
		14'b00100011001101:	sigmoid_prime = 18'b000000110001000011;
		14'b00100011001110:	sigmoid_prime = 18'b000000110000111101;
		14'b00100011001111:	sigmoid_prime = 18'b000000110000110111;
		14'b00100011010000:	sigmoid_prime = 18'b000000110000110001;
		14'b00100011010001:	sigmoid_prime = 18'b000000110000101011;
		14'b00100011010010:	sigmoid_prime = 18'b000000110000100101;
		14'b00100011010011:	sigmoid_prime = 18'b000000110000011111;
		14'b00100011010100:	sigmoid_prime = 18'b000000110000011010;
		14'b00100011010101:	sigmoid_prime = 18'b000000110000010100;
		14'b00100011010110:	sigmoid_prime = 18'b000000110000001110;
		14'b00100011010111:	sigmoid_prime = 18'b000000110000001000;
		14'b00100011011000:	sigmoid_prime = 18'b000000110000000010;
		14'b00100011011001:	sigmoid_prime = 18'b000000101111111100;
		14'b00100011011010:	sigmoid_prime = 18'b000000101111110110;
		14'b00100011011011:	sigmoid_prime = 18'b000000101111110000;
		14'b00100011011100:	sigmoid_prime = 18'b000000101111101011;
		14'b00100011011101:	sigmoid_prime = 18'b000000101111100101;
		14'b00100011011110:	sigmoid_prime = 18'b000000101111011111;
		14'b00100011011111:	sigmoid_prime = 18'b000000101111011001;
		14'b00100011100000:	sigmoid_prime = 18'b000000101111010011;
		14'b00100011100001:	sigmoid_prime = 18'b000000101111001110;
		14'b00100011100010:	sigmoid_prime = 18'b000000101111001000;
		14'b00100011100011:	sigmoid_prime = 18'b000000101111000010;
		14'b00100011100100:	sigmoid_prime = 18'b000000101110111100;
		14'b00100011100101:	sigmoid_prime = 18'b000000101110110111;
		14'b00100011100110:	sigmoid_prime = 18'b000000101110110001;
		14'b00100011100111:	sigmoid_prime = 18'b000000101110101011;
		14'b00100011101000:	sigmoid_prime = 18'b000000101110100110;
		14'b00100011101001:	sigmoid_prime = 18'b000000101110100000;
		14'b00100011101010:	sigmoid_prime = 18'b000000101110011010;
		14'b00100011101011:	sigmoid_prime = 18'b000000101110010101;
		14'b00100011101100:	sigmoid_prime = 18'b000000101110001111;
		14'b00100011101101:	sigmoid_prime = 18'b000000101110001001;
		14'b00100011101110:	sigmoid_prime = 18'b000000101110000100;
		14'b00100011101111:	sigmoid_prime = 18'b000000101101111110;
		14'b00100011110000:	sigmoid_prime = 18'b000000101101111000;
		14'b00100011110001:	sigmoid_prime = 18'b000000101101110011;
		14'b00100011110010:	sigmoid_prime = 18'b000000101101101101;
		14'b00100011110011:	sigmoid_prime = 18'b000000101101101000;
		14'b00100011110100:	sigmoid_prime = 18'b000000101101100010;
		14'b00100011110101:	sigmoid_prime = 18'b000000101101011100;
		14'b00100011110110:	sigmoid_prime = 18'b000000101101010111;
		14'b00100011110111:	sigmoid_prime = 18'b000000101101010001;
		14'b00100011111000:	sigmoid_prime = 18'b000000101101001100;
		14'b00100011111001:	sigmoid_prime = 18'b000000101101000110;
		14'b00100011111010:	sigmoid_prime = 18'b000000101101000001;
		14'b00100011111011:	sigmoid_prime = 18'b000000101100111011;
		14'b00100011111100:	sigmoid_prime = 18'b000000101100110110;
		14'b00100011111101:	sigmoid_prime = 18'b000000101100110000;
		14'b00100011111110:	sigmoid_prime = 18'b000000101100101011;
		14'b00100011111111:	sigmoid_prime = 18'b000000101100100101;
		14'b00100100000000:	sigmoid_prime = 18'b000000101100100000;
		14'b00100100000001:	sigmoid_prime = 18'b000000101100011011;
		14'b00100100000010:	sigmoid_prime = 18'b000000101100010101;
		14'b00100100000011:	sigmoid_prime = 18'b000000101100010000;
		14'b00100100000100:	sigmoid_prime = 18'b000000101100001010;
		14'b00100100000101:	sigmoid_prime = 18'b000000101100000101;
		14'b00100100000110:	sigmoid_prime = 18'b000000101100000000;
		14'b00100100000111:	sigmoid_prime = 18'b000000101011111010;
		14'b00100100001000:	sigmoid_prime = 18'b000000101011110101;
		14'b00100100001001:	sigmoid_prime = 18'b000000101011101111;
		14'b00100100001010:	sigmoid_prime = 18'b000000101011101010;
		14'b00100100001011:	sigmoid_prime = 18'b000000101011100101;
		14'b00100100001100:	sigmoid_prime = 18'b000000101011011111;
		14'b00100100001101:	sigmoid_prime = 18'b000000101011011010;
		14'b00100100001110:	sigmoid_prime = 18'b000000101011010101;
		14'b00100100001111:	sigmoid_prime = 18'b000000101011010000;
		14'b00100100010000:	sigmoid_prime = 18'b000000101011001010;
		14'b00100100010001:	sigmoid_prime = 18'b000000101011000101;
		14'b00100100010010:	sigmoid_prime = 18'b000000101011000000;
		14'b00100100010011:	sigmoid_prime = 18'b000000101010111010;
		14'b00100100010100:	sigmoid_prime = 18'b000000101010110101;
		14'b00100100010101:	sigmoid_prime = 18'b000000101010110000;
		14'b00100100010110:	sigmoid_prime = 18'b000000101010101011;
		14'b00100100010111:	sigmoid_prime = 18'b000000101010100110;
		14'b00100100011000:	sigmoid_prime = 18'b000000101010100000;
		14'b00100100011001:	sigmoid_prime = 18'b000000101010011011;
		14'b00100100011010:	sigmoid_prime = 18'b000000101010010110;
		14'b00100100011011:	sigmoid_prime = 18'b000000101010010001;
		14'b00100100011100:	sigmoid_prime = 18'b000000101010001100;
		14'b00100100011101:	sigmoid_prime = 18'b000000101010000110;
		14'b00100100011110:	sigmoid_prime = 18'b000000101010000001;
		14'b00100100011111:	sigmoid_prime = 18'b000000101001111100;
		14'b00100100100000:	sigmoid_prime = 18'b000000101001110111;
		14'b00100100100001:	sigmoid_prime = 18'b000000101001110010;
		14'b00100100100010:	sigmoid_prime = 18'b000000101001101101;
		14'b00100100100011:	sigmoid_prime = 18'b000000101001101000;
		14'b00100100100100:	sigmoid_prime = 18'b000000101001100011;
		14'b00100100100101:	sigmoid_prime = 18'b000000101001011101;
		14'b00100100100110:	sigmoid_prime = 18'b000000101001011000;
		14'b00100100100111:	sigmoid_prime = 18'b000000101001010011;
		14'b00100100101000:	sigmoid_prime = 18'b000000101001001110;
		14'b00100100101001:	sigmoid_prime = 18'b000000101001001001;
		14'b00100100101010:	sigmoid_prime = 18'b000000101001000100;
		14'b00100100101011:	sigmoid_prime = 18'b000000101000111111;
		14'b00100100101100:	sigmoid_prime = 18'b000000101000111010;
		14'b00100100101101:	sigmoid_prime = 18'b000000101000110101;
		14'b00100100101110:	sigmoid_prime = 18'b000000101000110000;
		14'b00100100101111:	sigmoid_prime = 18'b000000101000101011;
		14'b00100100110000:	sigmoid_prime = 18'b000000101000100110;
		14'b00100100110001:	sigmoid_prime = 18'b000000101000100001;
		14'b00100100110010:	sigmoid_prime = 18'b000000101000011100;
		14'b00100100110011:	sigmoid_prime = 18'b000000101000010111;
		14'b00100100110100:	sigmoid_prime = 18'b000000101000010010;
		14'b00100100110101:	sigmoid_prime = 18'b000000101000001101;
		14'b00100100110110:	sigmoid_prime = 18'b000000101000001001;
		14'b00100100110111:	sigmoid_prime = 18'b000000101000000100;
		14'b00100100111000:	sigmoid_prime = 18'b000000100111111111;
		14'b00100100111001:	sigmoid_prime = 18'b000000100111111010;
		14'b00100100111010:	sigmoid_prime = 18'b000000100111110101;
		14'b00100100111011:	sigmoid_prime = 18'b000000100111110000;
		14'b00100100111100:	sigmoid_prime = 18'b000000100111101011;
		14'b00100100111101:	sigmoid_prime = 18'b000000100111100110;
		14'b00100100111110:	sigmoid_prime = 18'b000000100111100001;
		14'b00100100111111:	sigmoid_prime = 18'b000000100111011101;
		14'b00100101000000:	sigmoid_prime = 18'b000000100111011000;
		14'b00100101000001:	sigmoid_prime = 18'b000000100111010011;
		14'b00100101000010:	sigmoid_prime = 18'b000000100111001110;
		14'b00100101000011:	sigmoid_prime = 18'b000000100111001001;
		14'b00100101000100:	sigmoid_prime = 18'b000000100111000101;
		14'b00100101000101:	sigmoid_prime = 18'b000000100111000000;
		14'b00100101000110:	sigmoid_prime = 18'b000000100110111011;
		14'b00100101000111:	sigmoid_prime = 18'b000000100110110110;
		14'b00100101001000:	sigmoid_prime = 18'b000000100110110001;
		14'b00100101001001:	sigmoid_prime = 18'b000000100110101101;
		14'b00100101001010:	sigmoid_prime = 18'b000000100110101000;
		14'b00100101001011:	sigmoid_prime = 18'b000000100110100011;
		14'b00100101001100:	sigmoid_prime = 18'b000000100110011111;
		14'b00100101001101:	sigmoid_prime = 18'b000000100110011010;
		14'b00100101001110:	sigmoid_prime = 18'b000000100110010101;
		14'b00100101001111:	sigmoid_prime = 18'b000000100110010000;
		14'b00100101010000:	sigmoid_prime = 18'b000000100110001100;
		14'b00100101010001:	sigmoid_prime = 18'b000000100110000111;
		14'b00100101010010:	sigmoid_prime = 18'b000000100110000010;
		14'b00100101010011:	sigmoid_prime = 18'b000000100101111110;
		14'b00100101010100:	sigmoid_prime = 18'b000000100101111001;
		14'b00100101010101:	sigmoid_prime = 18'b000000100101110100;
		14'b00100101010110:	sigmoid_prime = 18'b000000100101110000;
		14'b00100101010111:	sigmoid_prime = 18'b000000100101101011;
		14'b00100101011000:	sigmoid_prime = 18'b000000100101100111;
		14'b00100101011001:	sigmoid_prime = 18'b000000100101100010;
		14'b00100101011010:	sigmoid_prime = 18'b000000100101011101;
		14'b00100101011011:	sigmoid_prime = 18'b000000100101011001;
		14'b00100101011100:	sigmoid_prime = 18'b000000100101010100;
		14'b00100101011101:	sigmoid_prime = 18'b000000100101010000;
		14'b00100101011110:	sigmoid_prime = 18'b000000100101001011;
		14'b00100101011111:	sigmoid_prime = 18'b000000100101000110;
		14'b00100101100000:	sigmoid_prime = 18'b000000100101000010;
		14'b00100101100001:	sigmoid_prime = 18'b000000100100111101;
		14'b00100101100010:	sigmoid_prime = 18'b000000100100111001;
		14'b00100101100011:	sigmoid_prime = 18'b000000100100110100;
		14'b00100101100100:	sigmoid_prime = 18'b000000100100110000;
		14'b00100101100101:	sigmoid_prime = 18'b000000100100101011;
		14'b00100101100110:	sigmoid_prime = 18'b000000100100100111;
		14'b00100101100111:	sigmoid_prime = 18'b000000100100100010;
		14'b00100101101000:	sigmoid_prime = 18'b000000100100011110;
		14'b00100101101001:	sigmoid_prime = 18'b000000100100011001;
		14'b00100101101010:	sigmoid_prime = 18'b000000100100010101;
		14'b00100101101011:	sigmoid_prime = 18'b000000100100010000;
		14'b00100101101100:	sigmoid_prime = 18'b000000100100001100;
		14'b00100101101101:	sigmoid_prime = 18'b000000100100001000;
		14'b00100101101110:	sigmoid_prime = 18'b000000100100000011;
		14'b00100101101111:	sigmoid_prime = 18'b000000100011111111;
		14'b00100101110000:	sigmoid_prime = 18'b000000100011111010;
		14'b00100101110001:	sigmoid_prime = 18'b000000100011110110;
		14'b00100101110010:	sigmoid_prime = 18'b000000100011110001;
		14'b00100101110011:	sigmoid_prime = 18'b000000100011101101;
		14'b00100101110100:	sigmoid_prime = 18'b000000100011101001;
		14'b00100101110101:	sigmoid_prime = 18'b000000100011100100;
		14'b00100101110110:	sigmoid_prime = 18'b000000100011100000;
		14'b00100101110111:	sigmoid_prime = 18'b000000100011011100;
		14'b00100101111000:	sigmoid_prime = 18'b000000100011010111;
		14'b00100101111001:	sigmoid_prime = 18'b000000100011010011;
		14'b00100101111010:	sigmoid_prime = 18'b000000100011001111;
		14'b00100101111011:	sigmoid_prime = 18'b000000100011001010;
		14'b00100101111100:	sigmoid_prime = 18'b000000100011000110;
		14'b00100101111101:	sigmoid_prime = 18'b000000100011000010;
		14'b00100101111110:	sigmoid_prime = 18'b000000100010111101;
		14'b00100101111111:	sigmoid_prime = 18'b000000100010111001;
		14'b00100110000000:	sigmoid_prime = 18'b000000100010110101;
		14'b00100110000001:	sigmoid_prime = 18'b000000100010110000;
		14'b00100110000010:	sigmoid_prime = 18'b000000100010101100;
		14'b00100110000011:	sigmoid_prime = 18'b000000100010101000;
		14'b00100110000100:	sigmoid_prime = 18'b000000100010100100;
		14'b00100110000101:	sigmoid_prime = 18'b000000100010011111;
		14'b00100110000110:	sigmoid_prime = 18'b000000100010011011;
		14'b00100110000111:	sigmoid_prime = 18'b000000100010010111;
		14'b00100110001000:	sigmoid_prime = 18'b000000100010010011;
		14'b00100110001001:	sigmoid_prime = 18'b000000100010001111;
		14'b00100110001010:	sigmoid_prime = 18'b000000100010001010;
		14'b00100110001011:	sigmoid_prime = 18'b000000100010000110;
		14'b00100110001100:	sigmoid_prime = 18'b000000100010000010;
		14'b00100110001101:	sigmoid_prime = 18'b000000100001111110;
		14'b00100110001110:	sigmoid_prime = 18'b000000100001111010;
		14'b00100110001111:	sigmoid_prime = 18'b000000100001110101;
		14'b00100110010000:	sigmoid_prime = 18'b000000100001110001;
		14'b00100110010001:	sigmoid_prime = 18'b000000100001101101;
		14'b00100110010010:	sigmoid_prime = 18'b000000100001101001;
		14'b00100110010011:	sigmoid_prime = 18'b000000100001100101;
		14'b00100110010100:	sigmoid_prime = 18'b000000100001100001;
		14'b00100110010101:	sigmoid_prime = 18'b000000100001011101;
		14'b00100110010110:	sigmoid_prime = 18'b000000100001011001;
		14'b00100110010111:	sigmoid_prime = 18'b000000100001010100;
		14'b00100110011000:	sigmoid_prime = 18'b000000100001010000;
		14'b00100110011001:	sigmoid_prime = 18'b000000100001001100;
		14'b00100110011010:	sigmoid_prime = 18'b000000100001001000;
		14'b00100110011011:	sigmoid_prime = 18'b000000100001000100;
		14'b00100110011100:	sigmoid_prime = 18'b000000100001000000;
		14'b00100110011101:	sigmoid_prime = 18'b000000100000111100;
		14'b00100110011110:	sigmoid_prime = 18'b000000100000111000;
		14'b00100110011111:	sigmoid_prime = 18'b000000100000110100;
		14'b00100110100000:	sigmoid_prime = 18'b000000100000110000;
		14'b00100110100001:	sigmoid_prime = 18'b000000100000101100;
		14'b00100110100010:	sigmoid_prime = 18'b000000100000101000;
		14'b00100110100011:	sigmoid_prime = 18'b000000100000100100;
		14'b00100110100100:	sigmoid_prime = 18'b000000100000100000;
		14'b00100110100101:	sigmoid_prime = 18'b000000100000011100;
		14'b00100110100110:	sigmoid_prime = 18'b000000100000011000;
		14'b00100110100111:	sigmoid_prime = 18'b000000100000010100;
		14'b00100110101000:	sigmoid_prime = 18'b000000100000010000;
		14'b00100110101001:	sigmoid_prime = 18'b000000100000001100;
		14'b00100110101010:	sigmoid_prime = 18'b000000100000001000;
		14'b00100110101011:	sigmoid_prime = 18'b000000100000000100;
		14'b00100110101100:	sigmoid_prime = 18'b000000100000000000;
		14'b00100110101101:	sigmoid_prime = 18'b000000011111111100;
		14'b00100110101110:	sigmoid_prime = 18'b000000011111111000;
		14'b00100110101111:	sigmoid_prime = 18'b000000011111110100;
		14'b00100110110000:	sigmoid_prime = 18'b000000011111110000;
		14'b00100110110001:	sigmoid_prime = 18'b000000011111101100;
		14'b00100110110010:	sigmoid_prime = 18'b000000011111101001;
		14'b00100110110011:	sigmoid_prime = 18'b000000011111100101;
		14'b00100110110100:	sigmoid_prime = 18'b000000011111100001;
		14'b00100110110101:	sigmoid_prime = 18'b000000011111011101;
		14'b00100110110110:	sigmoid_prime = 18'b000000011111011001;
		14'b00100110110111:	sigmoid_prime = 18'b000000011111010101;
		14'b00100110111000:	sigmoid_prime = 18'b000000011111010001;
		14'b00100110111001:	sigmoid_prime = 18'b000000011111001101;
		14'b00100110111010:	sigmoid_prime = 18'b000000011111001010;
		14'b00100110111011:	sigmoid_prime = 18'b000000011111000110;
		14'b00100110111100:	sigmoid_prime = 18'b000000011111000010;
		14'b00100110111101:	sigmoid_prime = 18'b000000011110111110;
		14'b00100110111110:	sigmoid_prime = 18'b000000011110111010;
		14'b00100110111111:	sigmoid_prime = 18'b000000011110110111;
		14'b00100111000000:	sigmoid_prime = 18'b000000011110110011;
		14'b00100111000001:	sigmoid_prime = 18'b000000011110101111;
		14'b00100111000010:	sigmoid_prime = 18'b000000011110101011;
		14'b00100111000011:	sigmoid_prime = 18'b000000011110100111;
		14'b00100111000100:	sigmoid_prime = 18'b000000011110100100;
		14'b00100111000101:	sigmoid_prime = 18'b000000011110100000;
		14'b00100111000110:	sigmoid_prime = 18'b000000011110011100;
		14'b00100111000111:	sigmoid_prime = 18'b000000011110011000;
		14'b00100111001000:	sigmoid_prime = 18'b000000011110010101;
		14'b00100111001001:	sigmoid_prime = 18'b000000011110010001;
		14'b00100111001010:	sigmoid_prime = 18'b000000011110001101;
		14'b00100111001011:	sigmoid_prime = 18'b000000011110001001;
		14'b00100111001100:	sigmoid_prime = 18'b000000011110000110;
		14'b00100111001101:	sigmoid_prime = 18'b000000011110000010;
		14'b00100111001110:	sigmoid_prime = 18'b000000011101111110;
		14'b00100111001111:	sigmoid_prime = 18'b000000011101111011;
		14'b00100111010000:	sigmoid_prime = 18'b000000011101110111;
		14'b00100111010001:	sigmoid_prime = 18'b000000011101110011;
		14'b00100111010010:	sigmoid_prime = 18'b000000011101110000;
		14'b00100111010011:	sigmoid_prime = 18'b000000011101101100;
		14'b00100111010100:	sigmoid_prime = 18'b000000011101101000;
		14'b00100111010101:	sigmoid_prime = 18'b000000011101100101;
		14'b00100111010110:	sigmoid_prime = 18'b000000011101100001;
		14'b00100111010111:	sigmoid_prime = 18'b000000011101011101;
		14'b00100111011000:	sigmoid_prime = 18'b000000011101011010;
		14'b00100111011001:	sigmoid_prime = 18'b000000011101010110;
		14'b00100111011010:	sigmoid_prime = 18'b000000011101010011;
		14'b00100111011011:	sigmoid_prime = 18'b000000011101001111;
		14'b00100111011100:	sigmoid_prime = 18'b000000011101001011;
		14'b00100111011101:	sigmoid_prime = 18'b000000011101001000;
		14'b00100111011110:	sigmoid_prime = 18'b000000011101000100;
		14'b00100111011111:	sigmoid_prime = 18'b000000011101000001;
		14'b00100111100000:	sigmoid_prime = 18'b000000011100111101;
		14'b00100111100001:	sigmoid_prime = 18'b000000011100111001;
		14'b00100111100010:	sigmoid_prime = 18'b000000011100110110;
		14'b00100111100011:	sigmoid_prime = 18'b000000011100110010;
		14'b00100111100100:	sigmoid_prime = 18'b000000011100101111;
		14'b00100111100101:	sigmoid_prime = 18'b000000011100101011;
		14'b00100111100110:	sigmoid_prime = 18'b000000011100101000;
		14'b00100111100111:	sigmoid_prime = 18'b000000011100100100;
		14'b00100111101000:	sigmoid_prime = 18'b000000011100100001;
		14'b00100111101001:	sigmoid_prime = 18'b000000011100011101;
		14'b00100111101010:	sigmoid_prime = 18'b000000011100011010;
		14'b00100111101011:	sigmoid_prime = 18'b000000011100010110;
		14'b00100111101100:	sigmoid_prime = 18'b000000011100010011;
		14'b00100111101101:	sigmoid_prime = 18'b000000011100001111;
		14'b00100111101110:	sigmoid_prime = 18'b000000011100001100;
		14'b00100111101111:	sigmoid_prime = 18'b000000011100001000;
		14'b00100111110000:	sigmoid_prime = 18'b000000011100000101;
		14'b00100111110001:	sigmoid_prime = 18'b000000011100000001;
		14'b00100111110010:	sigmoid_prime = 18'b000000011011111110;
		14'b00100111110011:	sigmoid_prime = 18'b000000011011111010;
		14'b00100111110100:	sigmoid_prime = 18'b000000011011110111;
		14'b00100111110101:	sigmoid_prime = 18'b000000011011110100;
		14'b00100111110110:	sigmoid_prime = 18'b000000011011110000;
		14'b00100111110111:	sigmoid_prime = 18'b000000011011101101;
		14'b00100111111000:	sigmoid_prime = 18'b000000011011101001;
		14'b00100111111001:	sigmoid_prime = 18'b000000011011100110;
		14'b00100111111010:	sigmoid_prime = 18'b000000011011100011;
		14'b00100111111011:	sigmoid_prime = 18'b000000011011011111;
		14'b00100111111100:	sigmoid_prime = 18'b000000011011011100;
		14'b00100111111101:	sigmoid_prime = 18'b000000011011011000;
		14'b00100111111110:	sigmoid_prime = 18'b000000011011010101;
		14'b00100111111111:	sigmoid_prime = 18'b000000011011010010;
		14'b00101000000000:	sigmoid_prime = 18'b000000011011001110;
		14'b00101000000001:	sigmoid_prime = 18'b000000011011001011;
		14'b00101000000010:	sigmoid_prime = 18'b000000011011001000;
		14'b00101000000011:	sigmoid_prime = 18'b000000011011000100;
		14'b00101000000100:	sigmoid_prime = 18'b000000011011000001;
		14'b00101000000101:	sigmoid_prime = 18'b000000011010111110;
		14'b00101000000110:	sigmoid_prime = 18'b000000011010111010;
		14'b00101000000111:	sigmoid_prime = 18'b000000011010110111;
		14'b00101000001000:	sigmoid_prime = 18'b000000011010110100;
		14'b00101000001001:	sigmoid_prime = 18'b000000011010110000;
		14'b00101000001010:	sigmoid_prime = 18'b000000011010101101;
		14'b00101000001011:	sigmoid_prime = 18'b000000011010101010;
		14'b00101000001100:	sigmoid_prime = 18'b000000011010100110;
		14'b00101000001101:	sigmoid_prime = 18'b000000011010100011;
		14'b00101000001110:	sigmoid_prime = 18'b000000011010100000;
		14'b00101000001111:	sigmoid_prime = 18'b000000011010011101;
		14'b00101000010000:	sigmoid_prime = 18'b000000011010011001;
		14'b00101000010001:	sigmoid_prime = 18'b000000011010010110;
		14'b00101000010010:	sigmoid_prime = 18'b000000011010010011;
		14'b00101000010011:	sigmoid_prime = 18'b000000011010010000;
		14'b00101000010100:	sigmoid_prime = 18'b000000011010001100;
		14'b00101000010101:	sigmoid_prime = 18'b000000011010001001;
		14'b00101000010110:	sigmoid_prime = 18'b000000011010000110;
		14'b00101000010111:	sigmoid_prime = 18'b000000011010000011;
		14'b00101000011000:	sigmoid_prime = 18'b000000011001111111;
		14'b00101000011001:	sigmoid_prime = 18'b000000011001111100;
		14'b00101000011010:	sigmoid_prime = 18'b000000011001111001;
		14'b00101000011011:	sigmoid_prime = 18'b000000011001110110;
		14'b00101000011100:	sigmoid_prime = 18'b000000011001110011;
		14'b00101000011101:	sigmoid_prime = 18'b000000011001101111;
		14'b00101000011110:	sigmoid_prime = 18'b000000011001101100;
		14'b00101000011111:	sigmoid_prime = 18'b000000011001101001;
		14'b00101000100000:	sigmoid_prime = 18'b000000011001100110;
		14'b00101000100001:	sigmoid_prime = 18'b000000011001100011;
		14'b00101000100010:	sigmoid_prime = 18'b000000011001100000;
		14'b00101000100011:	sigmoid_prime = 18'b000000011001011101;
		14'b00101000100100:	sigmoid_prime = 18'b000000011001011001;
		14'b00101000100101:	sigmoid_prime = 18'b000000011001010110;
		14'b00101000100110:	sigmoid_prime = 18'b000000011001010011;
		14'b00101000100111:	sigmoid_prime = 18'b000000011001010000;
		14'b00101000101000:	sigmoid_prime = 18'b000000011001001101;
		14'b00101000101001:	sigmoid_prime = 18'b000000011001001010;
		14'b00101000101010:	sigmoid_prime = 18'b000000011001000111;
		14'b00101000101011:	sigmoid_prime = 18'b000000011001000100;
		14'b00101000101100:	sigmoid_prime = 18'b000000011001000000;
		14'b00101000101101:	sigmoid_prime = 18'b000000011000111101;
		14'b00101000101110:	sigmoid_prime = 18'b000000011000111010;
		14'b00101000101111:	sigmoid_prime = 18'b000000011000110111;
		14'b00101000110000:	sigmoid_prime = 18'b000000011000110100;
		14'b00101000110001:	sigmoid_prime = 18'b000000011000110001;
		14'b00101000110010:	sigmoid_prime = 18'b000000011000101110;
		14'b00101000110011:	sigmoid_prime = 18'b000000011000101011;
		14'b00101000110100:	sigmoid_prime = 18'b000000011000101000;
		14'b00101000110101:	sigmoid_prime = 18'b000000011000100101;
		14'b00101000110110:	sigmoid_prime = 18'b000000011000100010;
		14'b00101000110111:	sigmoid_prime = 18'b000000011000011111;
		14'b00101000111000:	sigmoid_prime = 18'b000000011000011100;
		14'b00101000111001:	sigmoid_prime = 18'b000000011000011001;
		14'b00101000111010:	sigmoid_prime = 18'b000000011000010110;
		14'b00101000111011:	sigmoid_prime = 18'b000000011000010011;
		14'b00101000111100:	sigmoid_prime = 18'b000000011000010000;
		14'b00101000111101:	sigmoid_prime = 18'b000000011000001101;
		14'b00101000111110:	sigmoid_prime = 18'b000000011000001010;
		14'b00101000111111:	sigmoid_prime = 18'b000000011000000111;
		14'b00101001000000:	sigmoid_prime = 18'b000000011000000100;
		14'b00101001000001:	sigmoid_prime = 18'b000000011000000001;
		14'b00101001000010:	sigmoid_prime = 18'b000000010111111110;
		14'b00101001000011:	sigmoid_prime = 18'b000000010111111011;
		14'b00101001000100:	sigmoid_prime = 18'b000000010111111000;
		14'b00101001000101:	sigmoid_prime = 18'b000000010111110101;
		14'b00101001000110:	sigmoid_prime = 18'b000000010111110010;
		14'b00101001000111:	sigmoid_prime = 18'b000000010111101111;
		14'b00101001001000:	sigmoid_prime = 18'b000000010111101100;
		14'b00101001001001:	sigmoid_prime = 18'b000000010111101001;
		14'b00101001001010:	sigmoid_prime = 18'b000000010111100110;
		14'b00101001001011:	sigmoid_prime = 18'b000000010111100100;
		14'b00101001001100:	sigmoid_prime = 18'b000000010111100001;
		14'b00101001001101:	sigmoid_prime = 18'b000000010111011110;
		14'b00101001001110:	sigmoid_prime = 18'b000000010111011011;
		14'b00101001001111:	sigmoid_prime = 18'b000000010111011000;
		14'b00101001010000:	sigmoid_prime = 18'b000000010111010101;
		14'b00101001010001:	sigmoid_prime = 18'b000000010111010010;
		14'b00101001010010:	sigmoid_prime = 18'b000000010111001111;
		14'b00101001010011:	sigmoid_prime = 18'b000000010111001100;
		14'b00101001010100:	sigmoid_prime = 18'b000000010111001010;
		14'b00101001010101:	sigmoid_prime = 18'b000000010111000111;
		14'b00101001010110:	sigmoid_prime = 18'b000000010111000100;
		14'b00101001010111:	sigmoid_prime = 18'b000000010111000001;
		14'b00101001011000:	sigmoid_prime = 18'b000000010110111110;
		14'b00101001011001:	sigmoid_prime = 18'b000000010110111011;
		14'b00101001011010:	sigmoid_prime = 18'b000000010110111000;
		14'b00101001011011:	sigmoid_prime = 18'b000000010110110110;
		14'b00101001011100:	sigmoid_prime = 18'b000000010110110011;
		14'b00101001011101:	sigmoid_prime = 18'b000000010110110000;
		14'b00101001011110:	sigmoid_prime = 18'b000000010110101101;
		14'b00101001011111:	sigmoid_prime = 18'b000000010110101010;
		14'b00101001100000:	sigmoid_prime = 18'b000000010110101000;
		14'b00101001100001:	sigmoid_prime = 18'b000000010110100101;
		14'b00101001100010:	sigmoid_prime = 18'b000000010110100010;
		14'b00101001100011:	sigmoid_prime = 18'b000000010110011111;
		14'b00101001100100:	sigmoid_prime = 18'b000000010110011100;
		14'b00101001100101:	sigmoid_prime = 18'b000000010110011010;
		14'b00101001100110:	sigmoid_prime = 18'b000000010110010111;
		14'b00101001100111:	sigmoid_prime = 18'b000000010110010100;
		14'b00101001101000:	sigmoid_prime = 18'b000000010110010001;
		14'b00101001101001:	sigmoid_prime = 18'b000000010110001111;
		14'b00101001101010:	sigmoid_prime = 18'b000000010110001100;
		14'b00101001101011:	sigmoid_prime = 18'b000000010110001001;
		14'b00101001101100:	sigmoid_prime = 18'b000000010110000110;
		14'b00101001101101:	sigmoid_prime = 18'b000000010110000100;
		14'b00101001101110:	sigmoid_prime = 18'b000000010110000001;
		14'b00101001101111:	sigmoid_prime = 18'b000000010101111110;
		14'b00101001110000:	sigmoid_prime = 18'b000000010101111100;
		14'b00101001110001:	sigmoid_prime = 18'b000000010101111001;
		14'b00101001110010:	sigmoid_prime = 18'b000000010101110110;
		14'b00101001110011:	sigmoid_prime = 18'b000000010101110011;
		14'b00101001110100:	sigmoid_prime = 18'b000000010101110001;
		14'b00101001110101:	sigmoid_prime = 18'b000000010101101110;
		14'b00101001110110:	sigmoid_prime = 18'b000000010101101011;
		14'b00101001110111:	sigmoid_prime = 18'b000000010101101001;
		14'b00101001111000:	sigmoid_prime = 18'b000000010101100110;
		14'b00101001111001:	sigmoid_prime = 18'b000000010101100011;
		14'b00101001111010:	sigmoid_prime = 18'b000000010101100001;
		14'b00101001111011:	sigmoid_prime = 18'b000000010101011110;
		14'b00101001111100:	sigmoid_prime = 18'b000000010101011011;
		14'b00101001111101:	sigmoid_prime = 18'b000000010101011001;
		14'b00101001111110:	sigmoid_prime = 18'b000000010101010110;
		14'b00101001111111:	sigmoid_prime = 18'b000000010101010011;
		14'b00101010000000:	sigmoid_prime = 18'b000000010101010001;
		14'b00101010000001:	sigmoid_prime = 18'b000000010101001110;
		14'b00101010000010:	sigmoid_prime = 18'b000000010101001100;
		14'b00101010000011:	sigmoid_prime = 18'b000000010101001001;
		14'b00101010000100:	sigmoid_prime = 18'b000000010101000110;
		14'b00101010000101:	sigmoid_prime = 18'b000000010101000100;
		14'b00101010000110:	sigmoid_prime = 18'b000000010101000001;
		14'b00101010000111:	sigmoid_prime = 18'b000000010100111110;
		14'b00101010001000:	sigmoid_prime = 18'b000000010100111100;
		14'b00101010001001:	sigmoid_prime = 18'b000000010100111001;
		14'b00101010001010:	sigmoid_prime = 18'b000000010100110111;
		14'b00101010001011:	sigmoid_prime = 18'b000000010100110100;
		14'b00101010001100:	sigmoid_prime = 18'b000000010100110010;
		14'b00101010001101:	sigmoid_prime = 18'b000000010100101111;
		14'b00101010001110:	sigmoid_prime = 18'b000000010100101100;
		14'b00101010001111:	sigmoid_prime = 18'b000000010100101010;
		14'b00101010010000:	sigmoid_prime = 18'b000000010100100111;
		14'b00101010010001:	sigmoid_prime = 18'b000000010100100101;
		14'b00101010010010:	sigmoid_prime = 18'b000000010100100010;
		14'b00101010010011:	sigmoid_prime = 18'b000000010100100000;
		14'b00101010010100:	sigmoid_prime = 18'b000000010100011101;
		14'b00101010010101:	sigmoid_prime = 18'b000000010100011011;
		14'b00101010010110:	sigmoid_prime = 18'b000000010100011000;
		14'b00101010010111:	sigmoid_prime = 18'b000000010100010110;
		14'b00101010011000:	sigmoid_prime = 18'b000000010100010011;
		14'b00101010011001:	sigmoid_prime = 18'b000000010100010001;
		14'b00101010011010:	sigmoid_prime = 18'b000000010100001110;
		14'b00101010011011:	sigmoid_prime = 18'b000000010100001100;
		14'b00101010011100:	sigmoid_prime = 18'b000000010100001001;
		14'b00101010011101:	sigmoid_prime = 18'b000000010100000111;
		14'b00101010011110:	sigmoid_prime = 18'b000000010100000100;
		14'b00101010011111:	sigmoid_prime = 18'b000000010100000010;
		14'b00101010100000:	sigmoid_prime = 18'b000000010011111111;
		14'b00101010100001:	sigmoid_prime = 18'b000000010011111101;
		14'b00101010100010:	sigmoid_prime = 18'b000000010011111010;
		14'b00101010100011:	sigmoid_prime = 18'b000000010011111000;
		14'b00101010100100:	sigmoid_prime = 18'b000000010011110101;
		14'b00101010100101:	sigmoid_prime = 18'b000000010011110011;
		14'b00101010100110:	sigmoid_prime = 18'b000000010011110000;
		14'b00101010100111:	sigmoid_prime = 18'b000000010011101110;
		14'b00101010101000:	sigmoid_prime = 18'b000000010011101011;
		14'b00101010101001:	sigmoid_prime = 18'b000000010011101001;
		14'b00101010101010:	sigmoid_prime = 18'b000000010011100111;
		14'b00101010101011:	sigmoid_prime = 18'b000000010011100100;
		14'b00101010101100:	sigmoid_prime = 18'b000000010011100010;
		14'b00101010101101:	sigmoid_prime = 18'b000000010011011111;
		14'b00101010101110:	sigmoid_prime = 18'b000000010011011101;
		14'b00101010101111:	sigmoid_prime = 18'b000000010011011011;
		14'b00101010110000:	sigmoid_prime = 18'b000000010011011000;
		14'b00101010110001:	sigmoid_prime = 18'b000000010011010110;
		14'b00101010110010:	sigmoid_prime = 18'b000000010011010011;
		14'b00101010110011:	sigmoid_prime = 18'b000000010011010001;
		14'b00101010110100:	sigmoid_prime = 18'b000000010011001111;
		14'b00101010110101:	sigmoid_prime = 18'b000000010011001100;
		14'b00101010110110:	sigmoid_prime = 18'b000000010011001010;
		14'b00101010110111:	sigmoid_prime = 18'b000000010011000111;
		14'b00101010111000:	sigmoid_prime = 18'b000000010011000101;
		14'b00101010111001:	sigmoid_prime = 18'b000000010011000011;
		14'b00101010111010:	sigmoid_prime = 18'b000000010011000000;
		14'b00101010111011:	sigmoid_prime = 18'b000000010010111110;
		14'b00101010111100:	sigmoid_prime = 18'b000000010010111100;
		14'b00101010111101:	sigmoid_prime = 18'b000000010010111001;
		14'b00101010111110:	sigmoid_prime = 18'b000000010010110111;
		14'b00101010111111:	sigmoid_prime = 18'b000000010010110101;
		14'b00101011000000:	sigmoid_prime = 18'b000000010010110010;
		14'b00101011000001:	sigmoid_prime = 18'b000000010010110000;
		14'b00101011000010:	sigmoid_prime = 18'b000000010010101110;
		14'b00101011000011:	sigmoid_prime = 18'b000000010010101011;
		14'b00101011000100:	sigmoid_prime = 18'b000000010010101001;
		14'b00101011000101:	sigmoid_prime = 18'b000000010010100111;
		14'b00101011000110:	sigmoid_prime = 18'b000000010010100100;
		14'b00101011000111:	sigmoid_prime = 18'b000000010010100010;
		14'b00101011001000:	sigmoid_prime = 18'b000000010010100000;
		14'b00101011001001:	sigmoid_prime = 18'b000000010010011110;
		14'b00101011001010:	sigmoid_prime = 18'b000000010010011011;
		14'b00101011001011:	sigmoid_prime = 18'b000000010010011001;
		14'b00101011001100:	sigmoid_prime = 18'b000000010010010111;
		14'b00101011001101:	sigmoid_prime = 18'b000000010010010100;
		14'b00101011001110:	sigmoid_prime = 18'b000000010010010010;
		14'b00101011001111:	sigmoid_prime = 18'b000000010010010000;
		14'b00101011010000:	sigmoid_prime = 18'b000000010010001110;
		14'b00101011010001:	sigmoid_prime = 18'b000000010010001011;
		14'b00101011010010:	sigmoid_prime = 18'b000000010010001001;
		14'b00101011010011:	sigmoid_prime = 18'b000000010010000111;
		14'b00101011010100:	sigmoid_prime = 18'b000000010010000101;
		14'b00101011010101:	sigmoid_prime = 18'b000000010010000010;
		14'b00101011010110:	sigmoid_prime = 18'b000000010010000000;
		14'b00101011010111:	sigmoid_prime = 18'b000000010001111110;
		14'b00101011011000:	sigmoid_prime = 18'b000000010001111100;
		14'b00101011011001:	sigmoid_prime = 18'b000000010001111001;
		14'b00101011011010:	sigmoid_prime = 18'b000000010001110111;
		14'b00101011011011:	sigmoid_prime = 18'b000000010001110101;
		14'b00101011011100:	sigmoid_prime = 18'b000000010001110011;
		14'b00101011011101:	sigmoid_prime = 18'b000000010001110001;
		14'b00101011011110:	sigmoid_prime = 18'b000000010001101110;
		14'b00101011011111:	sigmoid_prime = 18'b000000010001101100;
		14'b00101011100000:	sigmoid_prime = 18'b000000010001101010;
		14'b00101011100001:	sigmoid_prime = 18'b000000010001101000;
		14'b00101011100010:	sigmoid_prime = 18'b000000010001100110;
		14'b00101011100011:	sigmoid_prime = 18'b000000010001100100;
		14'b00101011100100:	sigmoid_prime = 18'b000000010001100001;
		14'b00101011100101:	sigmoid_prime = 18'b000000010001011111;
		14'b00101011100110:	sigmoid_prime = 18'b000000010001011101;
		14'b00101011100111:	sigmoid_prime = 18'b000000010001011011;
		14'b00101011101000:	sigmoid_prime = 18'b000000010001011001;
		14'b00101011101001:	sigmoid_prime = 18'b000000010001010111;
		14'b00101011101010:	sigmoid_prime = 18'b000000010001010100;
		14'b00101011101011:	sigmoid_prime = 18'b000000010001010010;
		14'b00101011101100:	sigmoid_prime = 18'b000000010001010000;
		14'b00101011101101:	sigmoid_prime = 18'b000000010001001110;
		14'b00101011101110:	sigmoid_prime = 18'b000000010001001100;
		14'b00101011101111:	sigmoid_prime = 18'b000000010001001010;
		14'b00101011110000:	sigmoid_prime = 18'b000000010001001000;
		14'b00101011110001:	sigmoid_prime = 18'b000000010001000101;
		14'b00101011110010:	sigmoid_prime = 18'b000000010001000011;
		14'b00101011110011:	sigmoid_prime = 18'b000000010001000001;
		14'b00101011110100:	sigmoid_prime = 18'b000000010000111111;
		14'b00101011110101:	sigmoid_prime = 18'b000000010000111101;
		14'b00101011110110:	sigmoid_prime = 18'b000000010000111011;
		14'b00101011110111:	sigmoid_prime = 18'b000000010000111001;
		14'b00101011111000:	sigmoid_prime = 18'b000000010000110111;
		14'b00101011111001:	sigmoid_prime = 18'b000000010000110101;
		14'b00101011111010:	sigmoid_prime = 18'b000000010000110011;
		14'b00101011111011:	sigmoid_prime = 18'b000000010000110000;
		14'b00101011111100:	sigmoid_prime = 18'b000000010000101110;
		14'b00101011111101:	sigmoid_prime = 18'b000000010000101100;
		14'b00101011111110:	sigmoid_prime = 18'b000000010000101010;
		14'b00101011111111:	sigmoid_prime = 18'b000000010000101000;
		14'b00101100000000:	sigmoid_prime = 18'b000000010000100110;
		14'b00101100000001:	sigmoid_prime = 18'b000000010000100100;
		14'b00101100000010:	sigmoid_prime = 18'b000000010000100010;
		14'b00101100000011:	sigmoid_prime = 18'b000000010000100000;
		14'b00101100000100:	sigmoid_prime = 18'b000000010000011110;
		14'b00101100000101:	sigmoid_prime = 18'b000000010000011100;
		14'b00101100000110:	sigmoid_prime = 18'b000000010000011010;
		14'b00101100000111:	sigmoid_prime = 18'b000000010000011000;
		14'b00101100001000:	sigmoid_prime = 18'b000000010000010110;
		14'b00101100001001:	sigmoid_prime = 18'b000000010000010100;
		14'b00101100001010:	sigmoid_prime = 18'b000000010000010010;
		14'b00101100001011:	sigmoid_prime = 18'b000000010000010000;
		14'b00101100001100:	sigmoid_prime = 18'b000000010000001110;
		14'b00101100001101:	sigmoid_prime = 18'b000000010000001100;
		14'b00101100001110:	sigmoid_prime = 18'b000000010000001010;
		14'b00101100001111:	sigmoid_prime = 18'b000000010000001000;
		14'b00101100010000:	sigmoid_prime = 18'b000000010000000110;
		14'b00101100010001:	sigmoid_prime = 18'b000000010000000100;
		14'b00101100010010:	sigmoid_prime = 18'b000000010000000010;
		14'b00101100010011:	sigmoid_prime = 18'b000000010000000000;
		14'b00101100010100:	sigmoid_prime = 18'b000000001111111110;
		14'b00101100010101:	sigmoid_prime = 18'b000000001111111100;
		14'b00101100010110:	sigmoid_prime = 18'b000000001111111010;
		14'b00101100010111:	sigmoid_prime = 18'b000000001111111000;
		14'b00101100011000:	sigmoid_prime = 18'b000000001111110110;
		14'b00101100011001:	sigmoid_prime = 18'b000000001111110100;
		14'b00101100011010:	sigmoid_prime = 18'b000000001111110010;
		14'b00101100011011:	sigmoid_prime = 18'b000000001111110000;
		14'b00101100011100:	sigmoid_prime = 18'b000000001111101110;
		14'b00101100011101:	sigmoid_prime = 18'b000000001111101100;
		14'b00101100011110:	sigmoid_prime = 18'b000000001111101010;
		14'b00101100011111:	sigmoid_prime = 18'b000000001111101000;
		14'b00101100100000:	sigmoid_prime = 18'b000000001111100110;
		14'b00101100100001:	sigmoid_prime = 18'b000000001111100100;
		14'b00101100100010:	sigmoid_prime = 18'b000000001111100010;
		14'b00101100100011:	sigmoid_prime = 18'b000000001111100000;
		14'b00101100100100:	sigmoid_prime = 18'b000000001111011111;
		14'b00101100100101:	sigmoid_prime = 18'b000000001111011101;
		14'b00101100100110:	sigmoid_prime = 18'b000000001111011011;
		14'b00101100100111:	sigmoid_prime = 18'b000000001111011001;
		14'b00101100101000:	sigmoid_prime = 18'b000000001111010111;
		14'b00101100101001:	sigmoid_prime = 18'b000000001111010101;
		14'b00101100101010:	sigmoid_prime = 18'b000000001111010011;
		14'b00101100101011:	sigmoid_prime = 18'b000000001111010001;
		14'b00101100101100:	sigmoid_prime = 18'b000000001111001111;
		14'b00101100101101:	sigmoid_prime = 18'b000000001111001101;
		14'b00101100101110:	sigmoid_prime = 18'b000000001111001011;
		14'b00101100101111:	sigmoid_prime = 18'b000000001111001010;
		14'b00101100110000:	sigmoid_prime = 18'b000000001111001000;
		14'b00101100110001:	sigmoid_prime = 18'b000000001111000110;
		14'b00101100110010:	sigmoid_prime = 18'b000000001111000100;
		14'b00101100110011:	sigmoid_prime = 18'b000000001111000010;
		14'b00101100110100:	sigmoid_prime = 18'b000000001111000000;
		14'b00101100110101:	sigmoid_prime = 18'b000000001110111110;
		14'b00101100110110:	sigmoid_prime = 18'b000000001110111101;
		14'b00101100110111:	sigmoid_prime = 18'b000000001110111011;
		14'b00101100111000:	sigmoid_prime = 18'b000000001110111001;
		14'b00101100111001:	sigmoid_prime = 18'b000000001110110111;
		14'b00101100111010:	sigmoid_prime = 18'b000000001110110101;
		14'b00101100111011:	sigmoid_prime = 18'b000000001110110011;
		14'b00101100111100:	sigmoid_prime = 18'b000000001110110001;
		14'b00101100111101:	sigmoid_prime = 18'b000000001110110000;
		14'b00101100111110:	sigmoid_prime = 18'b000000001110101110;
		14'b00101100111111:	sigmoid_prime = 18'b000000001110101100;
		14'b00101101000000:	sigmoid_prime = 18'b000000001110101010;
		14'b00101101000001:	sigmoid_prime = 18'b000000001110101000;
		14'b00101101000010:	sigmoid_prime = 18'b000000001110100111;
		14'b00101101000011:	sigmoid_prime = 18'b000000001110100101;
		14'b00101101000100:	sigmoid_prime = 18'b000000001110100011;
		14'b00101101000101:	sigmoid_prime = 18'b000000001110100001;
		14'b00101101000110:	sigmoid_prime = 18'b000000001110011111;
		14'b00101101000111:	sigmoid_prime = 18'b000000001110011110;
		14'b00101101001000:	sigmoid_prime = 18'b000000001110011100;
		14'b00101101001001:	sigmoid_prime = 18'b000000001110011010;
		14'b00101101001010:	sigmoid_prime = 18'b000000001110011000;
		14'b00101101001011:	sigmoid_prime = 18'b000000001110010110;
		14'b00101101001100:	sigmoid_prime = 18'b000000001110010101;
		14'b00101101001101:	sigmoid_prime = 18'b000000001110010011;
		14'b00101101001110:	sigmoid_prime = 18'b000000001110010001;
		14'b00101101001111:	sigmoid_prime = 18'b000000001110001111;
		14'b00101101010000:	sigmoid_prime = 18'b000000001110001101;
		14'b00101101010001:	sigmoid_prime = 18'b000000001110001100;
		14'b00101101010010:	sigmoid_prime = 18'b000000001110001010;
		14'b00101101010011:	sigmoid_prime = 18'b000000001110001000;
		14'b00101101010100:	sigmoid_prime = 18'b000000001110000110;
		14'b00101101010101:	sigmoid_prime = 18'b000000001110000101;
		14'b00101101010110:	sigmoid_prime = 18'b000000001110000011;
		14'b00101101010111:	sigmoid_prime = 18'b000000001110000001;
		14'b00101101011000:	sigmoid_prime = 18'b000000001101111111;
		14'b00101101011001:	sigmoid_prime = 18'b000000001101111110;
		14'b00101101011010:	sigmoid_prime = 18'b000000001101111100;
		14'b00101101011011:	sigmoid_prime = 18'b000000001101111010;
		14'b00101101011100:	sigmoid_prime = 18'b000000001101111001;
		14'b00101101011101:	sigmoid_prime = 18'b000000001101110111;
		14'b00101101011110:	sigmoid_prime = 18'b000000001101110101;
		14'b00101101011111:	sigmoid_prime = 18'b000000001101110011;
		14'b00101101100000:	sigmoid_prime = 18'b000000001101110010;
		14'b00101101100001:	sigmoid_prime = 18'b000000001101110000;
		14'b00101101100010:	sigmoid_prime = 18'b000000001101101110;
		14'b00101101100011:	sigmoid_prime = 18'b000000001101101101;
		14'b00101101100100:	sigmoid_prime = 18'b000000001101101011;
		14'b00101101100101:	sigmoid_prime = 18'b000000001101101001;
		14'b00101101100110:	sigmoid_prime = 18'b000000001101100111;
		14'b00101101100111:	sigmoid_prime = 18'b000000001101100110;
		14'b00101101101000:	sigmoid_prime = 18'b000000001101100100;
		14'b00101101101001:	sigmoid_prime = 18'b000000001101100010;
		14'b00101101101010:	sigmoid_prime = 18'b000000001101100001;
		14'b00101101101011:	sigmoid_prime = 18'b000000001101011111;
		14'b00101101101100:	sigmoid_prime = 18'b000000001101011101;
		14'b00101101101101:	sigmoid_prime = 18'b000000001101011100;
		14'b00101101101110:	sigmoid_prime = 18'b000000001101011010;
		14'b00101101101111:	sigmoid_prime = 18'b000000001101011000;
		14'b00101101110000:	sigmoid_prime = 18'b000000001101010111;
		14'b00101101110001:	sigmoid_prime = 18'b000000001101010101;
		14'b00101101110010:	sigmoid_prime = 18'b000000001101010011;
		14'b00101101110011:	sigmoid_prime = 18'b000000001101010010;
		14'b00101101110100:	sigmoid_prime = 18'b000000001101010000;
		14'b00101101110101:	sigmoid_prime = 18'b000000001101001110;
		14'b00101101110110:	sigmoid_prime = 18'b000000001101001101;
		14'b00101101110111:	sigmoid_prime = 18'b000000001101001011;
		14'b00101101111000:	sigmoid_prime = 18'b000000001101001010;
		14'b00101101111001:	sigmoid_prime = 18'b000000001101001000;
		14'b00101101111010:	sigmoid_prime = 18'b000000001101000110;
		14'b00101101111011:	sigmoid_prime = 18'b000000001101000101;
		14'b00101101111100:	sigmoid_prime = 18'b000000001101000011;
		14'b00101101111101:	sigmoid_prime = 18'b000000001101000001;
		14'b00101101111110:	sigmoid_prime = 18'b000000001101000000;
		14'b00101101111111:	sigmoid_prime = 18'b000000001100111110;
		14'b00101110000000:	sigmoid_prime = 18'b000000001100111101;
		14'b00101110000001:	sigmoid_prime = 18'b000000001100111011;
		14'b00101110000010:	sigmoid_prime = 18'b000000001100111001;
		14'b00101110000011:	sigmoid_prime = 18'b000000001100111000;
		14'b00101110000100:	sigmoid_prime = 18'b000000001100110110;
		14'b00101110000101:	sigmoid_prime = 18'b000000001100110101;
		14'b00101110000110:	sigmoid_prime = 18'b000000001100110011;
		14'b00101110000111:	sigmoid_prime = 18'b000000001100110001;
		14'b00101110001000:	sigmoid_prime = 18'b000000001100110000;
		14'b00101110001001:	sigmoid_prime = 18'b000000001100101110;
		14'b00101110001010:	sigmoid_prime = 18'b000000001100101101;
		14'b00101110001011:	sigmoid_prime = 18'b000000001100101011;
		14'b00101110001100:	sigmoid_prime = 18'b000000001100101001;
		14'b00101110001101:	sigmoid_prime = 18'b000000001100101000;
		14'b00101110001110:	sigmoid_prime = 18'b000000001100100110;
		14'b00101110001111:	sigmoid_prime = 18'b000000001100100101;
		14'b00101110010000:	sigmoid_prime = 18'b000000001100100011;
		14'b00101110010001:	sigmoid_prime = 18'b000000001100100010;
		14'b00101110010010:	sigmoid_prime = 18'b000000001100100000;
		14'b00101110010011:	sigmoid_prime = 18'b000000001100011111;
		14'b00101110010100:	sigmoid_prime = 18'b000000001100011101;
		14'b00101110010101:	sigmoid_prime = 18'b000000001100011011;
		14'b00101110010110:	sigmoid_prime = 18'b000000001100011010;
		14'b00101110010111:	sigmoid_prime = 18'b000000001100011000;
		14'b00101110011000:	sigmoid_prime = 18'b000000001100010111;
		14'b00101110011001:	sigmoid_prime = 18'b000000001100010101;
		14'b00101110011010:	sigmoid_prime = 18'b000000001100010100;
		14'b00101110011011:	sigmoid_prime = 18'b000000001100010010;
		14'b00101110011100:	sigmoid_prime = 18'b000000001100010001;
		14'b00101110011101:	sigmoid_prime = 18'b000000001100001111;
		14'b00101110011110:	sigmoid_prime = 18'b000000001100001110;
		14'b00101110011111:	sigmoid_prime = 18'b000000001100001100;
		14'b00101110100000:	sigmoid_prime = 18'b000000001100001011;
		14'b00101110100001:	sigmoid_prime = 18'b000000001100001001;
		14'b00101110100010:	sigmoid_prime = 18'b000000001100001000;
		14'b00101110100011:	sigmoid_prime = 18'b000000001100000110;
		14'b00101110100100:	sigmoid_prime = 18'b000000001100000101;
		14'b00101110100101:	sigmoid_prime = 18'b000000001100000011;
		14'b00101110100110:	sigmoid_prime = 18'b000000001100000010;
		14'b00101110100111:	sigmoid_prime = 18'b000000001100000000;
		14'b00101110101000:	sigmoid_prime = 18'b000000001011111111;
		14'b00101110101001:	sigmoid_prime = 18'b000000001011111101;
		14'b00101110101010:	sigmoid_prime = 18'b000000001011111100;
		14'b00101110101011:	sigmoid_prime = 18'b000000001011111010;
		14'b00101110101100:	sigmoid_prime = 18'b000000001011111001;
		14'b00101110101101:	sigmoid_prime = 18'b000000001011110111;
		14'b00101110101110:	sigmoid_prime = 18'b000000001011110110;
		14'b00101110101111:	sigmoid_prime = 18'b000000001011110100;
		14'b00101110110000:	sigmoid_prime = 18'b000000001011110011;
		14'b00101110110001:	sigmoid_prime = 18'b000000001011110001;
		14'b00101110110010:	sigmoid_prime = 18'b000000001011110000;
		14'b00101110110011:	sigmoid_prime = 18'b000000001011101110;
		14'b00101110110100:	sigmoid_prime = 18'b000000001011101101;
		14'b00101110110101:	sigmoid_prime = 18'b000000001011101011;
		14'b00101110110110:	sigmoid_prime = 18'b000000001011101010;
		14'b00101110110111:	sigmoid_prime = 18'b000000001011101001;
		14'b00101110111000:	sigmoid_prime = 18'b000000001011100111;
		14'b00101110111001:	sigmoid_prime = 18'b000000001011100110;
		14'b00101110111010:	sigmoid_prime = 18'b000000001011100100;
		14'b00101110111011:	sigmoid_prime = 18'b000000001011100011;
		14'b00101110111100:	sigmoid_prime = 18'b000000001011100001;
		14'b00101110111101:	sigmoid_prime = 18'b000000001011100000;
		14'b00101110111110:	sigmoid_prime = 18'b000000001011011111;
		14'b00101110111111:	sigmoid_prime = 18'b000000001011011101;
		14'b00101111000000:	sigmoid_prime = 18'b000000001011011100;
		14'b00101111000001:	sigmoid_prime = 18'b000000001011011010;
		14'b00101111000010:	sigmoid_prime = 18'b000000001011011001;
		14'b00101111000011:	sigmoid_prime = 18'b000000001011010111;
		14'b00101111000100:	sigmoid_prime = 18'b000000001011010110;
		14'b00101111000101:	sigmoid_prime = 18'b000000001011010101;
		14'b00101111000110:	sigmoid_prime = 18'b000000001011010011;
		14'b00101111000111:	sigmoid_prime = 18'b000000001011010010;
		14'b00101111001000:	sigmoid_prime = 18'b000000001011010000;
		14'b00101111001001:	sigmoid_prime = 18'b000000001011001111;
		14'b00101111001010:	sigmoid_prime = 18'b000000001011001110;
		14'b00101111001011:	sigmoid_prime = 18'b000000001011001100;
		14'b00101111001100:	sigmoid_prime = 18'b000000001011001011;
		14'b00101111001101:	sigmoid_prime = 18'b000000001011001001;
		14'b00101111001110:	sigmoid_prime = 18'b000000001011001000;
		14'b00101111001111:	sigmoid_prime = 18'b000000001011000111;
		14'b00101111010000:	sigmoid_prime = 18'b000000001011000101;
		14'b00101111010001:	sigmoid_prime = 18'b000000001011000100;
		14'b00101111010010:	sigmoid_prime = 18'b000000001011000011;
		14'b00101111010011:	sigmoid_prime = 18'b000000001011000001;
		14'b00101111010100:	sigmoid_prime = 18'b000000001011000000;
		14'b00101111010101:	sigmoid_prime = 18'b000000001010111110;
		14'b00101111010110:	sigmoid_prime = 18'b000000001010111101;
		14'b00101111010111:	sigmoid_prime = 18'b000000001010111100;
		14'b00101111011000:	sigmoid_prime = 18'b000000001010111010;
		14'b00101111011001:	sigmoid_prime = 18'b000000001010111001;
		14'b00101111011010:	sigmoid_prime = 18'b000000001010111000;
		14'b00101111011011:	sigmoid_prime = 18'b000000001010110110;
		14'b00101111011100:	sigmoid_prime = 18'b000000001010110101;
		14'b00101111011101:	sigmoid_prime = 18'b000000001010110100;
		14'b00101111011110:	sigmoid_prime = 18'b000000001010110010;
		14'b00101111011111:	sigmoid_prime = 18'b000000001010110001;
		14'b00101111100000:	sigmoid_prime = 18'b000000001010110000;
		14'b00101111100001:	sigmoid_prime = 18'b000000001010101110;
		14'b00101111100010:	sigmoid_prime = 18'b000000001010101101;
		14'b00101111100011:	sigmoid_prime = 18'b000000001010101100;
		14'b00101111100100:	sigmoid_prime = 18'b000000001010101010;
		14'b00101111100101:	sigmoid_prime = 18'b000000001010101001;
		14'b00101111100110:	sigmoid_prime = 18'b000000001010101000;
		14'b00101111100111:	sigmoid_prime = 18'b000000001010100110;
		14'b00101111101000:	sigmoid_prime = 18'b000000001010100101;
		14'b00101111101001:	sigmoid_prime = 18'b000000001010100100;
		14'b00101111101010:	sigmoid_prime = 18'b000000001010100010;
		14'b00101111101011:	sigmoid_prime = 18'b000000001010100001;
		14'b00101111101100:	sigmoid_prime = 18'b000000001010100000;
		14'b00101111101101:	sigmoid_prime = 18'b000000001010011110;
		14'b00101111101110:	sigmoid_prime = 18'b000000001010011101;
		14'b00101111101111:	sigmoid_prime = 18'b000000001010011100;
		14'b00101111110000:	sigmoid_prime = 18'b000000001010011011;
		14'b00101111110001:	sigmoid_prime = 18'b000000001010011001;
		14'b00101111110010:	sigmoid_prime = 18'b000000001010011000;
		14'b00101111110011:	sigmoid_prime = 18'b000000001010010111;
		14'b00101111110100:	sigmoid_prime = 18'b000000001010010101;
		14'b00101111110101:	sigmoid_prime = 18'b000000001010010100;
		14'b00101111110110:	sigmoid_prime = 18'b000000001010010011;
		14'b00101111110111:	sigmoid_prime = 18'b000000001010010001;
		14'b00101111111000:	sigmoid_prime = 18'b000000001010010000;
		14'b00101111111001:	sigmoid_prime = 18'b000000001010001111;
		14'b00101111111010:	sigmoid_prime = 18'b000000001010001110;
		14'b00101111111011:	sigmoid_prime = 18'b000000001010001100;
		14'b00101111111100:	sigmoid_prime = 18'b000000001010001011;
		14'b00101111111101:	sigmoid_prime = 18'b000000001010001010;
		14'b00101111111110:	sigmoid_prime = 18'b000000001010001001;
		14'b00101111111111:	sigmoid_prime = 18'b000000001010000111;
		14'b00110000000000:	sigmoid_prime = 18'b000000001010000110;
		14'b00110000000001:	sigmoid_prime = 18'b000000001010000101;
		14'b00110000000010:	sigmoid_prime = 18'b000000001010000100;
		14'b00110000000011:	sigmoid_prime = 18'b000000001010000010;
		14'b00110000000100:	sigmoid_prime = 18'b000000001010000001;
		14'b00110000000101:	sigmoid_prime = 18'b000000001010000000;
		14'b00110000000110:	sigmoid_prime = 18'b000000001001111111;
		14'b00110000000111:	sigmoid_prime = 18'b000000001001111101;
		14'b00110000001000:	sigmoid_prime = 18'b000000001001111100;
		14'b00110000001001:	sigmoid_prime = 18'b000000001001111011;
		14'b00110000001010:	sigmoid_prime = 18'b000000001001111010;
		14'b00110000001011:	sigmoid_prime = 18'b000000001001111000;
		14'b00110000001100:	sigmoid_prime = 18'b000000001001110111;
		14'b00110000001101:	sigmoid_prime = 18'b000000001001110110;
		14'b00110000001110:	sigmoid_prime = 18'b000000001001110101;
		14'b00110000001111:	sigmoid_prime = 18'b000000001001110100;
		14'b00110000010000:	sigmoid_prime = 18'b000000001001110010;
		14'b00110000010001:	sigmoid_prime = 18'b000000001001110001;
		14'b00110000010010:	sigmoid_prime = 18'b000000001001110000;
		14'b00110000010011:	sigmoid_prime = 18'b000000001001101111;
		14'b00110000010100:	sigmoid_prime = 18'b000000001001101101;
		14'b00110000010101:	sigmoid_prime = 18'b000000001001101100;
		14'b00110000010110:	sigmoid_prime = 18'b000000001001101011;
		14'b00110000010111:	sigmoid_prime = 18'b000000001001101010;
		14'b00110000011000:	sigmoid_prime = 18'b000000001001101001;
		14'b00110000011001:	sigmoid_prime = 18'b000000001001100111;
		14'b00110000011010:	sigmoid_prime = 18'b000000001001100110;
		14'b00110000011011:	sigmoid_prime = 18'b000000001001100101;
		14'b00110000011100:	sigmoid_prime = 18'b000000001001100100;
		14'b00110000011101:	sigmoid_prime = 18'b000000001001100011;
		14'b00110000011110:	sigmoid_prime = 18'b000000001001100001;
		14'b00110000011111:	sigmoid_prime = 18'b000000001001100000;
		14'b00110000100000:	sigmoid_prime = 18'b000000001001011111;
		14'b00110000100001:	sigmoid_prime = 18'b000000001001011110;
		14'b00110000100010:	sigmoid_prime = 18'b000000001001011101;
		14'b00110000100011:	sigmoid_prime = 18'b000000001001011100;
		14'b00110000100100:	sigmoid_prime = 18'b000000001001011010;
		14'b00110000100101:	sigmoid_prime = 18'b000000001001011001;
		14'b00110000100110:	sigmoid_prime = 18'b000000001001011000;
		14'b00110000100111:	sigmoid_prime = 18'b000000001001010111;
		14'b00110000101000:	sigmoid_prime = 18'b000000001001010110;
		14'b00110000101001:	sigmoid_prime = 18'b000000001001010101;
		14'b00110000101010:	sigmoid_prime = 18'b000000001001010011;
		14'b00110000101011:	sigmoid_prime = 18'b000000001001010010;
		14'b00110000101100:	sigmoid_prime = 18'b000000001001010001;
		14'b00110000101101:	sigmoid_prime = 18'b000000001001010000;
		14'b00110000101110:	sigmoid_prime = 18'b000000001001001111;
		14'b00110000101111:	sigmoid_prime = 18'b000000001001001110;
		14'b00110000110000:	sigmoid_prime = 18'b000000001001001100;
		14'b00110000110001:	sigmoid_prime = 18'b000000001001001011;
		14'b00110000110010:	sigmoid_prime = 18'b000000001001001010;
		14'b00110000110011:	sigmoid_prime = 18'b000000001001001001;
		14'b00110000110100:	sigmoid_prime = 18'b000000001001001000;
		14'b00110000110101:	sigmoid_prime = 18'b000000001001000111;
		14'b00110000110110:	sigmoid_prime = 18'b000000001001000110;
		14'b00110000110111:	sigmoid_prime = 18'b000000001001000101;
		14'b00110000111000:	sigmoid_prime = 18'b000000001001000011;
		14'b00110000111001:	sigmoid_prime = 18'b000000001001000010;
		14'b00110000111010:	sigmoid_prime = 18'b000000001001000001;
		14'b00110000111011:	sigmoid_prime = 18'b000000001001000000;
		14'b00110000111100:	sigmoid_prime = 18'b000000001000111111;
		14'b00110000111101:	sigmoid_prime = 18'b000000001000111110;
		14'b00110000111110:	sigmoid_prime = 18'b000000001000111101;
		14'b00110000111111:	sigmoid_prime = 18'b000000001000111100;
		14'b00110001000000:	sigmoid_prime = 18'b000000001000111010;
		14'b00110001000001:	sigmoid_prime = 18'b000000001000111001;
		14'b00110001000010:	sigmoid_prime = 18'b000000001000111000;
		14'b00110001000011:	sigmoid_prime = 18'b000000001000110111;
		14'b00110001000100:	sigmoid_prime = 18'b000000001000110110;
		14'b00110001000101:	sigmoid_prime = 18'b000000001000110101;
		14'b00110001000110:	sigmoid_prime = 18'b000000001000110100;
		14'b00110001000111:	sigmoid_prime = 18'b000000001000110011;
		14'b00110001001000:	sigmoid_prime = 18'b000000001000110010;
		14'b00110001001001:	sigmoid_prime = 18'b000000001000110001;
		14'b00110001001010:	sigmoid_prime = 18'b000000001000101111;
		14'b00110001001011:	sigmoid_prime = 18'b000000001000101110;
		14'b00110001001100:	sigmoid_prime = 18'b000000001000101101;
		14'b00110001001101:	sigmoid_prime = 18'b000000001000101100;
		14'b00110001001110:	sigmoid_prime = 18'b000000001000101011;
		14'b00110001001111:	sigmoid_prime = 18'b000000001000101010;
		14'b00110001010000:	sigmoid_prime = 18'b000000001000101001;
		14'b00110001010001:	sigmoid_prime = 18'b000000001000101000;
		14'b00110001010010:	sigmoid_prime = 18'b000000001000100111;
		14'b00110001010011:	sigmoid_prime = 18'b000000001000100110;
		14'b00110001010100:	sigmoid_prime = 18'b000000001000100101;
		14'b00110001010101:	sigmoid_prime = 18'b000000001000100100;
		14'b00110001010110:	sigmoid_prime = 18'b000000001000100011;
		14'b00110001010111:	sigmoid_prime = 18'b000000001000100001;
		14'b00110001011000:	sigmoid_prime = 18'b000000001000100000;
		14'b00110001011001:	sigmoid_prime = 18'b000000001000011111;
		14'b00110001011010:	sigmoid_prime = 18'b000000001000011110;
		14'b00110001011011:	sigmoid_prime = 18'b000000001000011101;
		14'b00110001011100:	sigmoid_prime = 18'b000000001000011100;
		14'b00110001011101:	sigmoid_prime = 18'b000000001000011011;
		14'b00110001011110:	sigmoid_prime = 18'b000000001000011010;
		14'b00110001011111:	sigmoid_prime = 18'b000000001000011001;
		14'b00110001100000:	sigmoid_prime = 18'b000000001000011000;
		14'b00110001100001:	sigmoid_prime = 18'b000000001000010111;
		14'b00110001100010:	sigmoid_prime = 18'b000000001000010110;
		14'b00110001100011:	sigmoid_prime = 18'b000000001000010101;
		14'b00110001100100:	sigmoid_prime = 18'b000000001000010100;
		14'b00110001100101:	sigmoid_prime = 18'b000000001000010011;
		14'b00110001100110:	sigmoid_prime = 18'b000000001000010010;
		14'b00110001100111:	sigmoid_prime = 18'b000000001000010001;
		14'b00110001101000:	sigmoid_prime = 18'b000000001000010000;
		14'b00110001101001:	sigmoid_prime = 18'b000000001000001111;
		14'b00110001101010:	sigmoid_prime = 18'b000000001000001110;
		14'b00110001101011:	sigmoid_prime = 18'b000000001000001101;
		14'b00110001101100:	sigmoid_prime = 18'b000000001000001100;
		14'b00110001101101:	sigmoid_prime = 18'b000000001000001011;
		14'b00110001101110:	sigmoid_prime = 18'b000000001000001010;
		14'b00110001101111:	sigmoid_prime = 18'b000000001000001001;
		14'b00110001110000:	sigmoid_prime = 18'b000000001000001000;
		14'b00110001110001:	sigmoid_prime = 18'b000000001000000111;
		14'b00110001110010:	sigmoid_prime = 18'b000000001000000110;
		14'b00110001110011:	sigmoid_prime = 18'b000000001000000101;
		14'b00110001110100:	sigmoid_prime = 18'b000000001000000100;
		14'b00110001110101:	sigmoid_prime = 18'b000000001000000011;
		14'b00110001110110:	sigmoid_prime = 18'b000000001000000010;
		14'b00110001110111:	sigmoid_prime = 18'b000000001000000001;
		14'b00110001111000:	sigmoid_prime = 18'b000000001000000000;
		14'b00110001111001:	sigmoid_prime = 18'b000000000111111111;
		14'b00110001111010:	sigmoid_prime = 18'b000000000111111110;
		14'b00110001111011:	sigmoid_prime = 18'b000000000111111101;
		14'b00110001111100:	sigmoid_prime = 18'b000000000111111100;
		14'b00110001111101:	sigmoid_prime = 18'b000000000111111011;
		14'b00110001111110:	sigmoid_prime = 18'b000000000111111010;
		14'b00110001111111:	sigmoid_prime = 18'b000000000111111001;
		14'b00110010000000:	sigmoid_prime = 18'b000000000111111000;
		14'b00110010000001:	sigmoid_prime = 18'b000000000111110111;
		14'b00110010000010:	sigmoid_prime = 18'b000000000111110110;
		14'b00110010000011:	sigmoid_prime = 18'b000000000111110101;
		14'b00110010000100:	sigmoid_prime = 18'b000000000111110100;
		14'b00110010000101:	sigmoid_prime = 18'b000000000111110011;
		14'b00110010000110:	sigmoid_prime = 18'b000000000111110010;
		14'b00110010000111:	sigmoid_prime = 18'b000000000111110001;
		14'b00110010001000:	sigmoid_prime = 18'b000000000111110000;
		14'b00110010001001:	sigmoid_prime = 18'b000000000111101111;
		14'b00110010001010:	sigmoid_prime = 18'b000000000111101110;
		14'b00110010001011:	sigmoid_prime = 18'b000000000111101101;
		14'b00110010001100:	sigmoid_prime = 18'b000000000111101100;
		14'b00110010001101:	sigmoid_prime = 18'b000000000111101011;
		14'b00110010001110:	sigmoid_prime = 18'b000000000111101010;
		14'b00110010001111:	sigmoid_prime = 18'b000000000111101001;
		14'b00110010010000:	sigmoid_prime = 18'b000000000111101000;
		14'b00110010010001:	sigmoid_prime = 18'b000000000111100111;
		14'b00110010010010:	sigmoid_prime = 18'b000000000111100110;
		14'b00110010010011:	sigmoid_prime = 18'b000000000111100101;
		14'b00110010010100:	sigmoid_prime = 18'b000000000111100100;
		14'b00110010010101:	sigmoid_prime = 18'b000000000111100011;
		14'b00110010010110:	sigmoid_prime = 18'b000000000111100010;
		14'b00110010010111:	sigmoid_prime = 18'b000000000111100010;
		14'b00110010011000:	sigmoid_prime = 18'b000000000111100001;
		14'b00110010011001:	sigmoid_prime = 18'b000000000111100000;
		14'b00110010011010:	sigmoid_prime = 18'b000000000111011111;
		14'b00110010011011:	sigmoid_prime = 18'b000000000111011110;
		14'b00110010011100:	sigmoid_prime = 18'b000000000111011101;
		14'b00110010011101:	sigmoid_prime = 18'b000000000111011100;
		14'b00110010011110:	sigmoid_prime = 18'b000000000111011011;
		14'b00110010011111:	sigmoid_prime = 18'b000000000111011010;
		14'b00110010100000:	sigmoid_prime = 18'b000000000111011001;
		14'b00110010100001:	sigmoid_prime = 18'b000000000111011000;
		14'b00110010100010:	sigmoid_prime = 18'b000000000111010111;
		14'b00110010100011:	sigmoid_prime = 18'b000000000111010110;
		14'b00110010100100:	sigmoid_prime = 18'b000000000111010110;
		14'b00110010100101:	sigmoid_prime = 18'b000000000111010101;
		14'b00110010100110:	sigmoid_prime = 18'b000000000111010100;
		14'b00110010100111:	sigmoid_prime = 18'b000000000111010011;
		14'b00110010101000:	sigmoid_prime = 18'b000000000111010010;
		14'b00110010101001:	sigmoid_prime = 18'b000000000111010001;
		14'b00110010101010:	sigmoid_prime = 18'b000000000111010000;
		14'b00110010101011:	sigmoid_prime = 18'b000000000111001111;
		14'b00110010101100:	sigmoid_prime = 18'b000000000111001110;
		14'b00110010101101:	sigmoid_prime = 18'b000000000111001101;
		14'b00110010101110:	sigmoid_prime = 18'b000000000111001100;
		14'b00110010101111:	sigmoid_prime = 18'b000000000111001100;
		14'b00110010110000:	sigmoid_prime = 18'b000000000111001011;
		14'b00110010110001:	sigmoid_prime = 18'b000000000111001010;
		14'b00110010110010:	sigmoid_prime = 18'b000000000111001001;
		14'b00110010110011:	sigmoid_prime = 18'b000000000111001000;
		14'b00110010110100:	sigmoid_prime = 18'b000000000111000111;
		14'b00110010110101:	sigmoid_prime = 18'b000000000111000110;
		14'b00110010110110:	sigmoid_prime = 18'b000000000111000101;
		14'b00110010110111:	sigmoid_prime = 18'b000000000111000100;
		14'b00110010111000:	sigmoid_prime = 18'b000000000111000100;
		14'b00110010111001:	sigmoid_prime = 18'b000000000111000011;
		14'b00110010111010:	sigmoid_prime = 18'b000000000111000010;
		14'b00110010111011:	sigmoid_prime = 18'b000000000111000001;
		14'b00110010111100:	sigmoid_prime = 18'b000000000111000000;
		14'b00110010111101:	sigmoid_prime = 18'b000000000110111111;
		14'b00110010111110:	sigmoid_prime = 18'b000000000110111110;
		14'b00110010111111:	sigmoid_prime = 18'b000000000110111101;
		14'b00110011000000:	sigmoid_prime = 18'b000000000110111101;
		14'b00110011000001:	sigmoid_prime = 18'b000000000110111100;
		14'b00110011000010:	sigmoid_prime = 18'b000000000110111011;
		14'b00110011000011:	sigmoid_prime = 18'b000000000110111010;
		14'b00110011000100:	sigmoid_prime = 18'b000000000110111001;
		14'b00110011000101:	sigmoid_prime = 18'b000000000110111000;
		14'b00110011000110:	sigmoid_prime = 18'b000000000110110111;
		14'b00110011000111:	sigmoid_prime = 18'b000000000110110111;
		14'b00110011001000:	sigmoid_prime = 18'b000000000110110110;
		14'b00110011001001:	sigmoid_prime = 18'b000000000110110101;
		14'b00110011001010:	sigmoid_prime = 18'b000000000110110100;
		14'b00110011001011:	sigmoid_prime = 18'b000000000110110011;
		14'b00110011001100:	sigmoid_prime = 18'b000000000110110010;
		14'b00110011001101:	sigmoid_prime = 18'b000000000110110001;
		14'b00110011001110:	sigmoid_prime = 18'b000000000110110001;
		14'b00110011001111:	sigmoid_prime = 18'b000000000110110000;
		14'b00110011010000:	sigmoid_prime = 18'b000000000110101111;
		14'b00110011010001:	sigmoid_prime = 18'b000000000110101110;
		14'b00110011010010:	sigmoid_prime = 18'b000000000110101101;
		14'b00110011010011:	sigmoid_prime = 18'b000000000110101100;
		14'b00110011010100:	sigmoid_prime = 18'b000000000110101100;
		14'b00110011010101:	sigmoid_prime = 18'b000000000110101011;
		14'b00110011010110:	sigmoid_prime = 18'b000000000110101010;
		14'b00110011010111:	sigmoid_prime = 18'b000000000110101001;
		14'b00110011011000:	sigmoid_prime = 18'b000000000110101000;
		14'b00110011011001:	sigmoid_prime = 18'b000000000110100111;
		14'b00110011011010:	sigmoid_prime = 18'b000000000110100111;
		14'b00110011011011:	sigmoid_prime = 18'b000000000110100110;
		14'b00110011011100:	sigmoid_prime = 18'b000000000110100101;
		14'b00110011011101:	sigmoid_prime = 18'b000000000110100100;
		14'b00110011011110:	sigmoid_prime = 18'b000000000110100011;
		14'b00110011011111:	sigmoid_prime = 18'b000000000110100011;
		14'b00110011100000:	sigmoid_prime = 18'b000000000110100010;
		14'b00110011100001:	sigmoid_prime = 18'b000000000110100001;
		14'b00110011100010:	sigmoid_prime = 18'b000000000110100000;
		14'b00110011100011:	sigmoid_prime = 18'b000000000110011111;
		14'b00110011100100:	sigmoid_prime = 18'b000000000110011110;
		14'b00110011100101:	sigmoid_prime = 18'b000000000110011110;
		14'b00110011100110:	sigmoid_prime = 18'b000000000110011101;
		14'b00110011100111:	sigmoid_prime = 18'b000000000110011100;
		14'b00110011101000:	sigmoid_prime = 18'b000000000110011011;
		14'b00110011101001:	sigmoid_prime = 18'b000000000110011010;
		14'b00110011101010:	sigmoid_prime = 18'b000000000110011010;
		14'b00110011101011:	sigmoid_prime = 18'b000000000110011001;
		14'b00110011101100:	sigmoid_prime = 18'b000000000110011000;
		14'b00110011101101:	sigmoid_prime = 18'b000000000110010111;
		14'b00110011101110:	sigmoid_prime = 18'b000000000110010110;
		14'b00110011101111:	sigmoid_prime = 18'b000000000110010110;
		14'b00110011110000:	sigmoid_prime = 18'b000000000110010101;
		14'b00110011110001:	sigmoid_prime = 18'b000000000110010100;
		14'b00110011110010:	sigmoid_prime = 18'b000000000110010011;
		14'b00110011110011:	sigmoid_prime = 18'b000000000110010011;
		14'b00110011110100:	sigmoid_prime = 18'b000000000110010010;
		14'b00110011110101:	sigmoid_prime = 18'b000000000110010001;
		14'b00110011110110:	sigmoid_prime = 18'b000000000110010000;
		14'b00110011110111:	sigmoid_prime = 18'b000000000110001111;
		14'b00110011111000:	sigmoid_prime = 18'b000000000110001111;
		14'b00110011111001:	sigmoid_prime = 18'b000000000110001110;
		14'b00110011111010:	sigmoid_prime = 18'b000000000110001101;
		14'b00110011111011:	sigmoid_prime = 18'b000000000110001100;
		14'b00110011111100:	sigmoid_prime = 18'b000000000110001100;
		14'b00110011111101:	sigmoid_prime = 18'b000000000110001011;
		14'b00110011111110:	sigmoid_prime = 18'b000000000110001010;
		14'b00110011111111:	sigmoid_prime = 18'b000000000110001001;
		14'b00110100000000:	sigmoid_prime = 18'b000000000110001000;
		14'b00110100000001:	sigmoid_prime = 18'b000000000110001000;
		14'b00110100000010:	sigmoid_prime = 18'b000000000110000111;
		14'b00110100000011:	sigmoid_prime = 18'b000000000110000110;
		14'b00110100000100:	sigmoid_prime = 18'b000000000110000101;
		14'b00110100000101:	sigmoid_prime = 18'b000000000110000101;
		14'b00110100000110:	sigmoid_prime = 18'b000000000110000100;
		14'b00110100000111:	sigmoid_prime = 18'b000000000110000011;
		14'b00110100001000:	sigmoid_prime = 18'b000000000110000010;
		14'b00110100001001:	sigmoid_prime = 18'b000000000110000010;
		14'b00110100001010:	sigmoid_prime = 18'b000000000110000001;
		14'b00110100001011:	sigmoid_prime = 18'b000000000110000000;
		14'b00110100001100:	sigmoid_prime = 18'b000000000101111111;
		14'b00110100001101:	sigmoid_prime = 18'b000000000101111111;
		14'b00110100001110:	sigmoid_prime = 18'b000000000101111110;
		14'b00110100001111:	sigmoid_prime = 18'b000000000101111101;
		14'b00110100010000:	sigmoid_prime = 18'b000000000101111100;
		14'b00110100010001:	sigmoid_prime = 18'b000000000101111100;
		14'b00110100010010:	sigmoid_prime = 18'b000000000101111011;
		14'b00110100010011:	sigmoid_prime = 18'b000000000101111010;
		14'b00110100010100:	sigmoid_prime = 18'b000000000101111001;
		14'b00110100010101:	sigmoid_prime = 18'b000000000101111001;
		14'b00110100010110:	sigmoid_prime = 18'b000000000101111000;
		14'b00110100010111:	sigmoid_prime = 18'b000000000101110111;
		14'b00110100011000:	sigmoid_prime = 18'b000000000101110110;
		14'b00110100011001:	sigmoid_prime = 18'b000000000101110110;
		14'b00110100011010:	sigmoid_prime = 18'b000000000101110101;
		14'b00110100011011:	sigmoid_prime = 18'b000000000101110100;
		14'b00110100011100:	sigmoid_prime = 18'b000000000101110100;
		14'b00110100011101:	sigmoid_prime = 18'b000000000101110011;
		14'b00110100011110:	sigmoid_prime = 18'b000000000101110010;
		14'b00110100011111:	sigmoid_prime = 18'b000000000101110001;
		14'b00110100100000:	sigmoid_prime = 18'b000000000101110001;
		14'b00110100100001:	sigmoid_prime = 18'b000000000101110000;
		14'b00110100100010:	sigmoid_prime = 18'b000000000101101111;
		14'b00110100100011:	sigmoid_prime = 18'b000000000101101111;
		14'b00110100100100:	sigmoid_prime = 18'b000000000101101110;
		14'b00110100100101:	sigmoid_prime = 18'b000000000101101101;
		14'b00110100100110:	sigmoid_prime = 18'b000000000101101100;
		14'b00110100100111:	sigmoid_prime = 18'b000000000101101100;
		14'b00110100101000:	sigmoid_prime = 18'b000000000101101011;
		14'b00110100101001:	sigmoid_prime = 18'b000000000101101010;
		14'b00110100101010:	sigmoid_prime = 18'b000000000101101010;
		14'b00110100101011:	sigmoid_prime = 18'b000000000101101001;
		14'b00110100101100:	sigmoid_prime = 18'b000000000101101000;
		14'b00110100101101:	sigmoid_prime = 18'b000000000101100111;
		14'b00110100101110:	sigmoid_prime = 18'b000000000101100111;
		14'b00110100101111:	sigmoid_prime = 18'b000000000101100110;
		14'b00110100110000:	sigmoid_prime = 18'b000000000101100101;
		14'b00110100110001:	sigmoid_prime = 18'b000000000101100101;
		14'b00110100110010:	sigmoid_prime = 18'b000000000101100100;
		14'b00110100110011:	sigmoid_prime = 18'b000000000101100011;
		14'b00110100110100:	sigmoid_prime = 18'b000000000101100011;
		14'b00110100110101:	sigmoid_prime = 18'b000000000101100010;
		14'b00110100110110:	sigmoid_prime = 18'b000000000101100001;
		14'b00110100110111:	sigmoid_prime = 18'b000000000101100001;
		14'b00110100111000:	sigmoid_prime = 18'b000000000101100000;
		14'b00110100111001:	sigmoid_prime = 18'b000000000101011111;
		14'b00110100111010:	sigmoid_prime = 18'b000000000101011110;
		14'b00110100111011:	sigmoid_prime = 18'b000000000101011110;
		14'b00110100111100:	sigmoid_prime = 18'b000000000101011101;
		14'b00110100111101:	sigmoid_prime = 18'b000000000101011100;
		14'b00110100111110:	sigmoid_prime = 18'b000000000101011100;
		14'b00110100111111:	sigmoid_prime = 18'b000000000101011011;
		14'b00110101000000:	sigmoid_prime = 18'b000000000101011010;
		14'b00110101000001:	sigmoid_prime = 18'b000000000101011010;
		14'b00110101000010:	sigmoid_prime = 18'b000000000101011001;
		14'b00110101000011:	sigmoid_prime = 18'b000000000101011000;
		14'b00110101000100:	sigmoid_prime = 18'b000000000101011000;
		14'b00110101000101:	sigmoid_prime = 18'b000000000101010111;
		14'b00110101000110:	sigmoid_prime = 18'b000000000101010110;
		14'b00110101000111:	sigmoid_prime = 18'b000000000101010110;
		14'b00110101001000:	sigmoid_prime = 18'b000000000101010101;
		14'b00110101001001:	sigmoid_prime = 18'b000000000101010100;
		14'b00110101001010:	sigmoid_prime = 18'b000000000101010100;
		14'b00110101001011:	sigmoid_prime = 18'b000000000101010011;
		14'b00110101001100:	sigmoid_prime = 18'b000000000101010010;
		14'b00110101001101:	sigmoid_prime = 18'b000000000101010010;
		14'b00110101001110:	sigmoid_prime = 18'b000000000101010001;
		14'b00110101001111:	sigmoid_prime = 18'b000000000101010000;
		14'b00110101010000:	sigmoid_prime = 18'b000000000101010000;
		14'b00110101010001:	sigmoid_prime = 18'b000000000101001111;
		14'b00110101010010:	sigmoid_prime = 18'b000000000101001110;
		14'b00110101010011:	sigmoid_prime = 18'b000000000101001110;
		14'b00110101010100:	sigmoid_prime = 18'b000000000101001101;
		14'b00110101010101:	sigmoid_prime = 18'b000000000101001100;
		14'b00110101010110:	sigmoid_prime = 18'b000000000101001100;
		14'b00110101010111:	sigmoid_prime = 18'b000000000101001011;
		14'b00110101011000:	sigmoid_prime = 18'b000000000101001011;
		14'b00110101011001:	sigmoid_prime = 18'b000000000101001010;
		14'b00110101011010:	sigmoid_prime = 18'b000000000101001001;
		14'b00110101011011:	sigmoid_prime = 18'b000000000101001001;
		14'b00110101011100:	sigmoid_prime = 18'b000000000101001000;
		14'b00110101011101:	sigmoid_prime = 18'b000000000101000111;
		14'b00110101011110:	sigmoid_prime = 18'b000000000101000111;
		14'b00110101011111:	sigmoid_prime = 18'b000000000101000110;
		14'b00110101100000:	sigmoid_prime = 18'b000000000101000101;
		14'b00110101100001:	sigmoid_prime = 18'b000000000101000101;
		14'b00110101100010:	sigmoid_prime = 18'b000000000101000100;
		14'b00110101100011:	sigmoid_prime = 18'b000000000101000100;
		14'b00110101100100:	sigmoid_prime = 18'b000000000101000011;
		14'b00110101100101:	sigmoid_prime = 18'b000000000101000010;
		14'b00110101100110:	sigmoid_prime = 18'b000000000101000010;
		14'b00110101100111:	sigmoid_prime = 18'b000000000101000001;
		14'b00110101101000:	sigmoid_prime = 18'b000000000101000000;
		14'b00110101101001:	sigmoid_prime = 18'b000000000101000000;
		14'b00110101101010:	sigmoid_prime = 18'b000000000100111111;
		14'b00110101101011:	sigmoid_prime = 18'b000000000100111111;
		14'b00110101101100:	sigmoid_prime = 18'b000000000100111110;
		14'b00110101101101:	sigmoid_prime = 18'b000000000100111101;
		14'b00110101101110:	sigmoid_prime = 18'b000000000100111101;
		14'b00110101101111:	sigmoid_prime = 18'b000000000100111100;
		14'b00110101110000:	sigmoid_prime = 18'b000000000100111011;
		14'b00110101110001:	sigmoid_prime = 18'b000000000100111011;
		14'b00110101110010:	sigmoid_prime = 18'b000000000100111010;
		14'b00110101110011:	sigmoid_prime = 18'b000000000100111010;
		14'b00110101110100:	sigmoid_prime = 18'b000000000100111001;
		14'b00110101110101:	sigmoid_prime = 18'b000000000100111000;
		14'b00110101110110:	sigmoid_prime = 18'b000000000100111000;
		14'b00110101110111:	sigmoid_prime = 18'b000000000100110111;
		14'b00110101111000:	sigmoid_prime = 18'b000000000100110111;
		14'b00110101111001:	sigmoid_prime = 18'b000000000100110110;
		14'b00110101111010:	sigmoid_prime = 18'b000000000100110101;
		14'b00110101111011:	sigmoid_prime = 18'b000000000100110101;
		14'b00110101111100:	sigmoid_prime = 18'b000000000100110100;
		14'b00110101111101:	sigmoid_prime = 18'b000000000100110100;
		14'b00110101111110:	sigmoid_prime = 18'b000000000100110011;
		14'b00110101111111:	sigmoid_prime = 18'b000000000100110010;
		14'b00110110000000:	sigmoid_prime = 18'b000000000100110010;
		14'b00110110000001:	sigmoid_prime = 18'b000000000100110001;
		14'b00110110000010:	sigmoid_prime = 18'b000000000100110001;
		14'b00110110000011:	sigmoid_prime = 18'b000000000100110000;
		14'b00110110000100:	sigmoid_prime = 18'b000000000100101111;
		14'b00110110000101:	sigmoid_prime = 18'b000000000100101111;
		14'b00110110000110:	sigmoid_prime = 18'b000000000100101110;
		14'b00110110000111:	sigmoid_prime = 18'b000000000100101110;
		14'b00110110001000:	sigmoid_prime = 18'b000000000100101101;
		14'b00110110001001:	sigmoid_prime = 18'b000000000100101100;
		14'b00110110001010:	sigmoid_prime = 18'b000000000100101100;
		14'b00110110001011:	sigmoid_prime = 18'b000000000100101011;
		14'b00110110001100:	sigmoid_prime = 18'b000000000100101011;
		14'b00110110001101:	sigmoid_prime = 18'b000000000100101010;
		14'b00110110001110:	sigmoid_prime = 18'b000000000100101001;
		14'b00110110001111:	sigmoid_prime = 18'b000000000100101001;
		14'b00110110010000:	sigmoid_prime = 18'b000000000100101000;
		14'b00110110010001:	sigmoid_prime = 18'b000000000100101000;
		14'b00110110010010:	sigmoid_prime = 18'b000000000100100111;
		14'b00110110010011:	sigmoid_prime = 18'b000000000100100111;
		14'b00110110010100:	sigmoid_prime = 18'b000000000100100110;
		14'b00110110010101:	sigmoid_prime = 18'b000000000100100101;
		14'b00110110010110:	sigmoid_prime = 18'b000000000100100101;
		14'b00110110010111:	sigmoid_prime = 18'b000000000100100100;
		14'b00110110011000:	sigmoid_prime = 18'b000000000100100100;
		14'b00110110011001:	sigmoid_prime = 18'b000000000100100011;
		14'b00110110011010:	sigmoid_prime = 18'b000000000100100011;
		14'b00110110011011:	sigmoid_prime = 18'b000000000100100010;
		14'b00110110011100:	sigmoid_prime = 18'b000000000100100001;
		14'b00110110011101:	sigmoid_prime = 18'b000000000100100001;
		14'b00110110011110:	sigmoid_prime = 18'b000000000100100000;
		14'b00110110011111:	sigmoid_prime = 18'b000000000100100000;
		14'b00110110100000:	sigmoid_prime = 18'b000000000100011111;
		14'b00110110100001:	sigmoid_prime = 18'b000000000100011111;
		14'b00110110100010:	sigmoid_prime = 18'b000000000100011110;
		14'b00110110100011:	sigmoid_prime = 18'b000000000100011110;
		14'b00110110100100:	sigmoid_prime = 18'b000000000100011101;
		14'b00110110100101:	sigmoid_prime = 18'b000000000100011100;
		14'b00110110100110:	sigmoid_prime = 18'b000000000100011100;
		14'b00110110100111:	sigmoid_prime = 18'b000000000100011011;
		14'b00110110101000:	sigmoid_prime = 18'b000000000100011011;
		14'b00110110101001:	sigmoid_prime = 18'b000000000100011010;
		14'b00110110101010:	sigmoid_prime = 18'b000000000100011010;
		14'b00110110101011:	sigmoid_prime = 18'b000000000100011001;
		14'b00110110101100:	sigmoid_prime = 18'b000000000100011001;
		14'b00110110101101:	sigmoid_prime = 18'b000000000100011000;
		14'b00110110101110:	sigmoid_prime = 18'b000000000100010111;
		14'b00110110101111:	sigmoid_prime = 18'b000000000100010111;
		14'b00110110110000:	sigmoid_prime = 18'b000000000100010110;
		14'b00110110110001:	sigmoid_prime = 18'b000000000100010110;
		14'b00110110110010:	sigmoid_prime = 18'b000000000100010101;
		14'b00110110110011:	sigmoid_prime = 18'b000000000100010101;
		14'b00110110110100:	sigmoid_prime = 18'b000000000100010100;
		14'b00110110110101:	sigmoid_prime = 18'b000000000100010100;
		14'b00110110110110:	sigmoid_prime = 18'b000000000100010011;
		14'b00110110110111:	sigmoid_prime = 18'b000000000100010011;
		14'b00110110111000:	sigmoid_prime = 18'b000000000100010010;
		14'b00110110111001:	sigmoid_prime = 18'b000000000100010010;
		14'b00110110111010:	sigmoid_prime = 18'b000000000100010001;
		14'b00110110111011:	sigmoid_prime = 18'b000000000100010000;
		14'b00110110111100:	sigmoid_prime = 18'b000000000100010000;
		14'b00110110111101:	sigmoid_prime = 18'b000000000100001111;
		14'b00110110111110:	sigmoid_prime = 18'b000000000100001111;
		14'b00110110111111:	sigmoid_prime = 18'b000000000100001110;
		14'b00110111000000:	sigmoid_prime = 18'b000000000100001110;
		14'b00110111000001:	sigmoid_prime = 18'b000000000100001101;
		14'b00110111000010:	sigmoid_prime = 18'b000000000100001101;
		14'b00110111000011:	sigmoid_prime = 18'b000000000100001100;
		14'b00110111000100:	sigmoid_prime = 18'b000000000100001100;
		14'b00110111000101:	sigmoid_prime = 18'b000000000100001011;
		14'b00110111000110:	sigmoid_prime = 18'b000000000100001011;
		14'b00110111000111:	sigmoid_prime = 18'b000000000100001010;
		14'b00110111001000:	sigmoid_prime = 18'b000000000100001010;
		14'b00110111001001:	sigmoid_prime = 18'b000000000100001001;
		14'b00110111001010:	sigmoid_prime = 18'b000000000100001001;
		14'b00110111001011:	sigmoid_prime = 18'b000000000100001000;
		14'b00110111001100:	sigmoid_prime = 18'b000000000100001000;
		14'b00110111001101:	sigmoid_prime = 18'b000000000100000111;
		14'b00110111001110:	sigmoid_prime = 18'b000000000100000111;
		14'b00110111001111:	sigmoid_prime = 18'b000000000100000110;
		14'b00110111010000:	sigmoid_prime = 18'b000000000100000110;
		14'b00110111010001:	sigmoid_prime = 18'b000000000100000101;
		14'b00110111010010:	sigmoid_prime = 18'b000000000100000100;
		14'b00110111010011:	sigmoid_prime = 18'b000000000100000100;
		14'b00110111010100:	sigmoid_prime = 18'b000000000100000011;
		14'b00110111010101:	sigmoid_prime = 18'b000000000100000011;
		14'b00110111010110:	sigmoid_prime = 18'b000000000100000010;
		14'b00110111010111:	sigmoid_prime = 18'b000000000100000010;
		14'b00110111011000:	sigmoid_prime = 18'b000000000100000001;
		14'b00110111011001:	sigmoid_prime = 18'b000000000100000001;
		14'b00110111011010:	sigmoid_prime = 18'b000000000100000000;
		14'b00110111011011:	sigmoid_prime = 18'b000000000100000000;
		14'b00110111011100:	sigmoid_prime = 18'b000000000011111111;
		14'b00110111011101:	sigmoid_prime = 18'b000000000011111111;
		14'b00110111011110:	sigmoid_prime = 18'b000000000011111110;
		14'b00110111011111:	sigmoid_prime = 18'b000000000011111110;
		14'b00110111100000:	sigmoid_prime = 18'b000000000011111101;
		14'b00110111100001:	sigmoid_prime = 18'b000000000011111101;
		14'b00110111100010:	sigmoid_prime = 18'b000000000011111100;
		14'b00110111100011:	sigmoid_prime = 18'b000000000011111100;
		14'b00110111100100:	sigmoid_prime = 18'b000000000011111011;
		14'b00110111100101:	sigmoid_prime = 18'b000000000011111011;
		14'b00110111100110:	sigmoid_prime = 18'b000000000011111011;
		14'b00110111100111:	sigmoid_prime = 18'b000000000011111010;
		14'b00110111101000:	sigmoid_prime = 18'b000000000011111010;
		14'b00110111101001:	sigmoid_prime = 18'b000000000011111001;
		14'b00110111101010:	sigmoid_prime = 18'b000000000011111001;
		14'b00110111101011:	sigmoid_prime = 18'b000000000011111000;
		14'b00110111101100:	sigmoid_prime = 18'b000000000011111000;
		14'b00110111101101:	sigmoid_prime = 18'b000000000011110111;
		14'b00110111101110:	sigmoid_prime = 18'b000000000011110111;
		14'b00110111101111:	sigmoid_prime = 18'b000000000011110110;
		14'b00110111110000:	sigmoid_prime = 18'b000000000011110110;
		14'b00110111110001:	sigmoid_prime = 18'b000000000011110101;
		14'b00110111110010:	sigmoid_prime = 18'b000000000011110101;
		14'b00110111110011:	sigmoid_prime = 18'b000000000011110100;
		14'b00110111110100:	sigmoid_prime = 18'b000000000011110100;
		14'b00110111110101:	sigmoid_prime = 18'b000000000011110011;
		14'b00110111110110:	sigmoid_prime = 18'b000000000011110011;
		14'b00110111110111:	sigmoid_prime = 18'b000000000011110010;
		14'b00110111111000:	sigmoid_prime = 18'b000000000011110010;
		14'b00110111111001:	sigmoid_prime = 18'b000000000011110001;
		14'b00110111111010:	sigmoid_prime = 18'b000000000011110001;
		14'b00110111111011:	sigmoid_prime = 18'b000000000011110000;
		14'b00110111111100:	sigmoid_prime = 18'b000000000011110000;
		14'b00110111111101:	sigmoid_prime = 18'b000000000011110000;
		14'b00110111111110:	sigmoid_prime = 18'b000000000011101111;
		14'b00110111111111:	sigmoid_prime = 18'b000000000011101111;
		14'b00111000000000:	sigmoid_prime = 18'b000000000011101110;
		14'b00111000000001:	sigmoid_prime = 18'b000000000011101110;
		14'b00111000000010:	sigmoid_prime = 18'b000000000011101101;
		14'b00111000000011:	sigmoid_prime = 18'b000000000011101101;
		14'b00111000000100:	sigmoid_prime = 18'b000000000011101100;
		14'b00111000000101:	sigmoid_prime = 18'b000000000011101100;
		14'b00111000000110:	sigmoid_prime = 18'b000000000011101011;
		14'b00111000000111:	sigmoid_prime = 18'b000000000011101011;
		14'b00111000001000:	sigmoid_prime = 18'b000000000011101010;
		14'b00111000001001:	sigmoid_prime = 18'b000000000011101010;
		14'b00111000001010:	sigmoid_prime = 18'b000000000011101010;
		14'b00111000001011:	sigmoid_prime = 18'b000000000011101001;
		14'b00111000001100:	sigmoid_prime = 18'b000000000011101001;
		14'b00111000001101:	sigmoid_prime = 18'b000000000011101000;
		14'b00111000001110:	sigmoid_prime = 18'b000000000011101000;
		14'b00111000001111:	sigmoid_prime = 18'b000000000011100111;
		14'b00111000010000:	sigmoid_prime = 18'b000000000011100111;
		14'b00111000010001:	sigmoid_prime = 18'b000000000011100110;
		14'b00111000010010:	sigmoid_prime = 18'b000000000011100110;
		14'b00111000010011:	sigmoid_prime = 18'b000000000011100101;
		14'b00111000010100:	sigmoid_prime = 18'b000000000011100101;
		14'b00111000010101:	sigmoid_prime = 18'b000000000011100101;
		14'b00111000010110:	sigmoid_prime = 18'b000000000011100100;
		14'b00111000010111:	sigmoid_prime = 18'b000000000011100100;
		14'b00111000011000:	sigmoid_prime = 18'b000000000011100011;
		14'b00111000011001:	sigmoid_prime = 18'b000000000011100011;
		14'b00111000011010:	sigmoid_prime = 18'b000000000011100010;
		14'b00111000011011:	sigmoid_prime = 18'b000000000011100010;
		14'b00111000011100:	sigmoid_prime = 18'b000000000011100001;
		14'b00111000011101:	sigmoid_prime = 18'b000000000011100001;
		14'b00111000011110:	sigmoid_prime = 18'b000000000011100001;
		14'b00111000011111:	sigmoid_prime = 18'b000000000011100000;
		14'b00111000100000:	sigmoid_prime = 18'b000000000011100000;
		14'b00111000100001:	sigmoid_prime = 18'b000000000011011111;
		14'b00111000100010:	sigmoid_prime = 18'b000000000011011111;
		14'b00111000100011:	sigmoid_prime = 18'b000000000011011110;
		14'b00111000100100:	sigmoid_prime = 18'b000000000011011110;
		14'b00111000100101:	sigmoid_prime = 18'b000000000011011110;
		14'b00111000100110:	sigmoid_prime = 18'b000000000011011101;
		14'b00111000100111:	sigmoid_prime = 18'b000000000011011101;
		14'b00111000101000:	sigmoid_prime = 18'b000000000011011100;
		14'b00111000101001:	sigmoid_prime = 18'b000000000011011100;
		14'b00111000101010:	sigmoid_prime = 18'b000000000011011011;
		14'b00111000101011:	sigmoid_prime = 18'b000000000011011011;
		14'b00111000101100:	sigmoid_prime = 18'b000000000011011010;
		14'b00111000101101:	sigmoid_prime = 18'b000000000011011010;
		14'b00111000101110:	sigmoid_prime = 18'b000000000011011010;
		14'b00111000101111:	sigmoid_prime = 18'b000000000011011001;
		14'b00111000110000:	sigmoid_prime = 18'b000000000011011001;
		14'b00111000110001:	sigmoid_prime = 18'b000000000011011000;
		14'b00111000110010:	sigmoid_prime = 18'b000000000011011000;
		14'b00111000110011:	sigmoid_prime = 18'b000000000011011000;
		14'b00111000110100:	sigmoid_prime = 18'b000000000011010111;
		14'b00111000110101:	sigmoid_prime = 18'b000000000011010111;
		14'b00111000110110:	sigmoid_prime = 18'b000000000011010110;
		14'b00111000110111:	sigmoid_prime = 18'b000000000011010110;
		14'b00111000111000:	sigmoid_prime = 18'b000000000011010101;
		14'b00111000111001:	sigmoid_prime = 18'b000000000011010101;
		14'b00111000111010:	sigmoid_prime = 18'b000000000011010101;
		14'b00111000111011:	sigmoid_prime = 18'b000000000011010100;
		14'b00111000111100:	sigmoid_prime = 18'b000000000011010100;
		14'b00111000111101:	sigmoid_prime = 18'b000000000011010011;
		14'b00111000111110:	sigmoid_prime = 18'b000000000011010011;
		14'b00111000111111:	sigmoid_prime = 18'b000000000011010011;
		14'b00111001000000:	sigmoid_prime = 18'b000000000011010010;
		14'b00111001000001:	sigmoid_prime = 18'b000000000011010010;
		14'b00111001000010:	sigmoid_prime = 18'b000000000011010001;
		14'b00111001000011:	sigmoid_prime = 18'b000000000011010001;
		14'b00111001000100:	sigmoid_prime = 18'b000000000011010000;
		14'b00111001000101:	sigmoid_prime = 18'b000000000011010000;
		14'b00111001000110:	sigmoid_prime = 18'b000000000011010000;
		14'b00111001000111:	sigmoid_prime = 18'b000000000011001111;
		14'b00111001001000:	sigmoid_prime = 18'b000000000011001111;
		14'b00111001001001:	sigmoid_prime = 18'b000000000011001110;
		14'b00111001001010:	sigmoid_prime = 18'b000000000011001110;
		14'b00111001001011:	sigmoid_prime = 18'b000000000011001110;
		14'b00111001001100:	sigmoid_prime = 18'b000000000011001101;
		14'b00111001001101:	sigmoid_prime = 18'b000000000011001101;
		14'b00111001001110:	sigmoid_prime = 18'b000000000011001100;
		14'b00111001001111:	sigmoid_prime = 18'b000000000011001100;
		14'b00111001010000:	sigmoid_prime = 18'b000000000011001100;
		14'b00111001010001:	sigmoid_prime = 18'b000000000011001011;
		14'b00111001010010:	sigmoid_prime = 18'b000000000011001011;
		14'b00111001010011:	sigmoid_prime = 18'b000000000011001010;
		14'b00111001010100:	sigmoid_prime = 18'b000000000011001010;
		14'b00111001010101:	sigmoid_prime = 18'b000000000011001010;
		14'b00111001010110:	sigmoid_prime = 18'b000000000011001001;
		14'b00111001010111:	sigmoid_prime = 18'b000000000011001001;
		14'b00111001011000:	sigmoid_prime = 18'b000000000011001000;
		14'b00111001011001:	sigmoid_prime = 18'b000000000011001000;
		14'b00111001011010:	sigmoid_prime = 18'b000000000011001000;
		14'b00111001011011:	sigmoid_prime = 18'b000000000011000111;
		14'b00111001011100:	sigmoid_prime = 18'b000000000011000111;
		14'b00111001011101:	sigmoid_prime = 18'b000000000011000111;
		14'b00111001011110:	sigmoid_prime = 18'b000000000011000110;
		14'b00111001011111:	sigmoid_prime = 18'b000000000011000110;
		14'b00111001100000:	sigmoid_prime = 18'b000000000011000101;
		14'b00111001100001:	sigmoid_prime = 18'b000000000011000101;
		14'b00111001100010:	sigmoid_prime = 18'b000000000011000101;
		14'b00111001100011:	sigmoid_prime = 18'b000000000011000100;
		14'b00111001100100:	sigmoid_prime = 18'b000000000011000100;
		14'b00111001100101:	sigmoid_prime = 18'b000000000011000011;
		14'b00111001100110:	sigmoid_prime = 18'b000000000011000011;
		14'b00111001100111:	sigmoid_prime = 18'b000000000011000011;
		14'b00111001101000:	sigmoid_prime = 18'b000000000011000010;
		14'b00111001101001:	sigmoid_prime = 18'b000000000011000010;
		14'b00111001101010:	sigmoid_prime = 18'b000000000011000010;
		14'b00111001101011:	sigmoid_prime = 18'b000000000011000001;
		14'b00111001101100:	sigmoid_prime = 18'b000000000011000001;
		14'b00111001101101:	sigmoid_prime = 18'b000000000011000000;
		14'b00111001101110:	sigmoid_prime = 18'b000000000011000000;
		14'b00111001101111:	sigmoid_prime = 18'b000000000011000000;
		14'b00111001110000:	sigmoid_prime = 18'b000000000010111111;
		14'b00111001110001:	sigmoid_prime = 18'b000000000010111111;
		14'b00111001110010:	sigmoid_prime = 18'b000000000010111111;
		14'b00111001110011:	sigmoid_prime = 18'b000000000010111110;
		14'b00111001110100:	sigmoid_prime = 18'b000000000010111110;
		14'b00111001110101:	sigmoid_prime = 18'b000000000010111101;
		14'b00111001110110:	sigmoid_prime = 18'b000000000010111101;
		14'b00111001110111:	sigmoid_prime = 18'b000000000010111101;
		14'b00111001111000:	sigmoid_prime = 18'b000000000010111100;
		14'b00111001111001:	sigmoid_prime = 18'b000000000010111100;
		14'b00111001111010:	sigmoid_prime = 18'b000000000010111100;
		14'b00111001111011:	sigmoid_prime = 18'b000000000010111011;
		14'b00111001111100:	sigmoid_prime = 18'b000000000010111011;
		14'b00111001111101:	sigmoid_prime = 18'b000000000010111010;
		14'b00111001111110:	sigmoid_prime = 18'b000000000010111010;
		14'b00111001111111:	sigmoid_prime = 18'b000000000010111010;
		14'b00111010000000:	sigmoid_prime = 18'b000000000010111001;
		14'b00111010000001:	sigmoid_prime = 18'b000000000010111001;
		14'b00111010000010:	sigmoid_prime = 18'b000000000010111001;
		14'b00111010000011:	sigmoid_prime = 18'b000000000010111000;
		14'b00111010000100:	sigmoid_prime = 18'b000000000010111000;
		14'b00111010000101:	sigmoid_prime = 18'b000000000010111000;
		14'b00111010000110:	sigmoid_prime = 18'b000000000010110111;
		14'b00111010000111:	sigmoid_prime = 18'b000000000010110111;
		14'b00111010001000:	sigmoid_prime = 18'b000000000010110111;
		14'b00111010001001:	sigmoid_prime = 18'b000000000010110110;
		14'b00111010001010:	sigmoid_prime = 18'b000000000010110110;
		14'b00111010001011:	sigmoid_prime = 18'b000000000010110101;
		14'b00111010001100:	sigmoid_prime = 18'b000000000010110101;
		14'b00111010001101:	sigmoid_prime = 18'b000000000010110101;
		14'b00111010001110:	sigmoid_prime = 18'b000000000010110100;
		14'b00111010001111:	sigmoid_prime = 18'b000000000010110100;
		14'b00111010010000:	sigmoid_prime = 18'b000000000010110100;
		14'b00111010010001:	sigmoid_prime = 18'b000000000010110011;
		14'b00111010010010:	sigmoid_prime = 18'b000000000010110011;
		14'b00111010010011:	sigmoid_prime = 18'b000000000010110011;
		14'b00111010010100:	sigmoid_prime = 18'b000000000010110010;
		14'b00111010010101:	sigmoid_prime = 18'b000000000010110010;
		14'b00111010010110:	sigmoid_prime = 18'b000000000010110010;
		14'b00111010010111:	sigmoid_prime = 18'b000000000010110001;
		14'b00111010011000:	sigmoid_prime = 18'b000000000010110001;
		14'b00111010011001:	sigmoid_prime = 18'b000000000010110001;
		14'b00111010011010:	sigmoid_prime = 18'b000000000010110000;
		14'b00111010011011:	sigmoid_prime = 18'b000000000010110000;
		14'b00111010011100:	sigmoid_prime = 18'b000000000010110000;
		14'b00111010011101:	sigmoid_prime = 18'b000000000010101111;
		14'b00111010011110:	sigmoid_prime = 18'b000000000010101111;
		14'b00111010011111:	sigmoid_prime = 18'b000000000010101110;
		14'b00111010100000:	sigmoid_prime = 18'b000000000010101110;
		14'b00111010100001:	sigmoid_prime = 18'b000000000010101110;
		14'b00111010100010:	sigmoid_prime = 18'b000000000010101101;
		14'b00111010100011:	sigmoid_prime = 18'b000000000010101101;
		14'b00111010100100:	sigmoid_prime = 18'b000000000010101101;
		14'b00111010100101:	sigmoid_prime = 18'b000000000010101100;
		14'b00111010100110:	sigmoid_prime = 18'b000000000010101100;
		14'b00111010100111:	sigmoid_prime = 18'b000000000010101100;
		14'b00111010101000:	sigmoid_prime = 18'b000000000010101011;
		14'b00111010101001:	sigmoid_prime = 18'b000000000010101011;
		14'b00111010101010:	sigmoid_prime = 18'b000000000010101011;
		14'b00111010101011:	sigmoid_prime = 18'b000000000010101010;
		14'b00111010101100:	sigmoid_prime = 18'b000000000010101010;
		14'b00111010101101:	sigmoid_prime = 18'b000000000010101010;
		14'b00111010101110:	sigmoid_prime = 18'b000000000010101001;
		14'b00111010101111:	sigmoid_prime = 18'b000000000010101001;
		14'b00111010110000:	sigmoid_prime = 18'b000000000010101001;
		14'b00111010110001:	sigmoid_prime = 18'b000000000010101000;
		14'b00111010110010:	sigmoid_prime = 18'b000000000010101000;
		14'b00111010110011:	sigmoid_prime = 18'b000000000010101000;
		14'b00111010110100:	sigmoid_prime = 18'b000000000010100111;
		14'b00111010110101:	sigmoid_prime = 18'b000000000010100111;
		14'b00111010110110:	sigmoid_prime = 18'b000000000010100111;
		14'b00111010110111:	sigmoid_prime = 18'b000000000010100110;
		14'b00111010111000:	sigmoid_prime = 18'b000000000010100110;
		14'b00111010111001:	sigmoid_prime = 18'b000000000010100110;
		14'b00111010111010:	sigmoid_prime = 18'b000000000010100110;
		14'b00111010111011:	sigmoid_prime = 18'b000000000010100101;
		14'b00111010111100:	sigmoid_prime = 18'b000000000010100101;
		14'b00111010111101:	sigmoid_prime = 18'b000000000010100101;
		14'b00111010111110:	sigmoid_prime = 18'b000000000010100100;
		14'b00111010111111:	sigmoid_prime = 18'b000000000010100100;
		14'b00111011000000:	sigmoid_prime = 18'b000000000010100100;
		14'b00111011000001:	sigmoid_prime = 18'b000000000010100011;
		14'b00111011000010:	sigmoid_prime = 18'b000000000010100011;
		14'b00111011000011:	sigmoid_prime = 18'b000000000010100011;
		14'b00111011000100:	sigmoid_prime = 18'b000000000010100010;
		14'b00111011000101:	sigmoid_prime = 18'b000000000010100010;
		14'b00111011000110:	sigmoid_prime = 18'b000000000010100010;
		14'b00111011000111:	sigmoid_prime = 18'b000000000010100001;
		14'b00111011001000:	sigmoid_prime = 18'b000000000010100001;
		14'b00111011001001:	sigmoid_prime = 18'b000000000010100001;
		14'b00111011001010:	sigmoid_prime = 18'b000000000010100000;
		14'b00111011001011:	sigmoid_prime = 18'b000000000010100000;
		14'b00111011001100:	sigmoid_prime = 18'b000000000010100000;
		14'b00111011001101:	sigmoid_prime = 18'b000000000010011111;
		14'b00111011001110:	sigmoid_prime = 18'b000000000010011111;
		14'b00111011001111:	sigmoid_prime = 18'b000000000010011111;
		14'b00111011010000:	sigmoid_prime = 18'b000000000010011111;
		14'b00111011010001:	sigmoid_prime = 18'b000000000010011110;
		14'b00111011010010:	sigmoid_prime = 18'b000000000010011110;
		14'b00111011010011:	sigmoid_prime = 18'b000000000010011110;
		14'b00111011010100:	sigmoid_prime = 18'b000000000010011101;
		14'b00111011010101:	sigmoid_prime = 18'b000000000010011101;
		14'b00111011010110:	sigmoid_prime = 18'b000000000010011101;
		14'b00111011010111:	sigmoid_prime = 18'b000000000010011100;
		14'b00111011011000:	sigmoid_prime = 18'b000000000010011100;
		14'b00111011011001:	sigmoid_prime = 18'b000000000010011100;
		14'b00111011011010:	sigmoid_prime = 18'b000000000010011011;
		14'b00111011011011:	sigmoid_prime = 18'b000000000010011011;
		14'b00111011011100:	sigmoid_prime = 18'b000000000010011011;
		14'b00111011011101:	sigmoid_prime = 18'b000000000010011011;
		14'b00111011011110:	sigmoid_prime = 18'b000000000010011010;
		14'b00111011011111:	sigmoid_prime = 18'b000000000010011010;
		14'b00111011100000:	sigmoid_prime = 18'b000000000010011010;
		14'b00111011100001:	sigmoid_prime = 18'b000000000010011001;
		14'b00111011100010:	sigmoid_prime = 18'b000000000010011001;
		14'b00111011100011:	sigmoid_prime = 18'b000000000010011001;
		14'b00111011100100:	sigmoid_prime = 18'b000000000010011000;
		14'b00111011100101:	sigmoid_prime = 18'b000000000010011000;
		14'b00111011100110:	sigmoid_prime = 18'b000000000010011000;
		14'b00111011100111:	sigmoid_prime = 18'b000000000010011000;
		14'b00111011101000:	sigmoid_prime = 18'b000000000010010111;
		14'b00111011101001:	sigmoid_prime = 18'b000000000010010111;
		14'b00111011101010:	sigmoid_prime = 18'b000000000010010111;
		14'b00111011101011:	sigmoid_prime = 18'b000000000010010110;
		14'b00111011101100:	sigmoid_prime = 18'b000000000010010110;
		14'b00111011101101:	sigmoid_prime = 18'b000000000010010110;
		14'b00111011101110:	sigmoid_prime = 18'b000000000010010110;
		14'b00111011101111:	sigmoid_prime = 18'b000000000010010101;
		14'b00111011110000:	sigmoid_prime = 18'b000000000010010101;
		14'b00111011110001:	sigmoid_prime = 18'b000000000010010101;
		14'b00111011110010:	sigmoid_prime = 18'b000000000010010100;
		14'b00111011110011:	sigmoid_prime = 18'b000000000010010100;
		14'b00111011110100:	sigmoid_prime = 18'b000000000010010100;
		14'b00111011110101:	sigmoid_prime = 18'b000000000010010011;
		14'b00111011110110:	sigmoid_prime = 18'b000000000010010011;
		14'b00111011110111:	sigmoid_prime = 18'b000000000010010011;
		14'b00111011111000:	sigmoid_prime = 18'b000000000010010011;
		14'b00111011111001:	sigmoid_prime = 18'b000000000010010010;
		14'b00111011111010:	sigmoid_prime = 18'b000000000010010010;
		14'b00111011111011:	sigmoid_prime = 18'b000000000010010010;
		14'b00111011111100:	sigmoid_prime = 18'b000000000010010001;
		14'b00111011111101:	sigmoid_prime = 18'b000000000010010001;
		14'b00111011111110:	sigmoid_prime = 18'b000000000010010001;
		14'b00111011111111:	sigmoid_prime = 18'b000000000010010001;
		14'b00111100000000:	sigmoid_prime = 18'b000000000010010000;
		14'b00111100000001:	sigmoid_prime = 18'b000000000010010000;
		14'b00111100000010:	sigmoid_prime = 18'b000000000010010000;
		14'b00111100000011:	sigmoid_prime = 18'b000000000010001111;
		14'b00111100000100:	sigmoid_prime = 18'b000000000010001111;
		14'b00111100000101:	sigmoid_prime = 18'b000000000010001111;
		14'b00111100000110:	sigmoid_prime = 18'b000000000010001111;
		14'b00111100000111:	sigmoid_prime = 18'b000000000010001110;
		14'b00111100001000:	sigmoid_prime = 18'b000000000010001110;
		14'b00111100001001:	sigmoid_prime = 18'b000000000010001110;
		14'b00111100001010:	sigmoid_prime = 18'b000000000010001110;
		14'b00111100001011:	sigmoid_prime = 18'b000000000010001101;
		14'b00111100001100:	sigmoid_prime = 18'b000000000010001101;
		14'b00111100001101:	sigmoid_prime = 18'b000000000010001101;
		14'b00111100001110:	sigmoid_prime = 18'b000000000010001100;
		14'b00111100001111:	sigmoid_prime = 18'b000000000010001100;
		14'b00111100010000:	sigmoid_prime = 18'b000000000010001100;
		14'b00111100010001:	sigmoid_prime = 18'b000000000010001100;
		14'b00111100010010:	sigmoid_prime = 18'b000000000010001011;
		14'b00111100010011:	sigmoid_prime = 18'b000000000010001011;
		14'b00111100010100:	sigmoid_prime = 18'b000000000010001011;
		14'b00111100010101:	sigmoid_prime = 18'b000000000010001011;
		14'b00111100010110:	sigmoid_prime = 18'b000000000010001010;
		14'b00111100010111:	sigmoid_prime = 18'b000000000010001010;
		14'b00111100011000:	sigmoid_prime = 18'b000000000010001010;
		14'b00111100011001:	sigmoid_prime = 18'b000000000010001001;
		14'b00111100011010:	sigmoid_prime = 18'b000000000010001001;
		14'b00111100011011:	sigmoid_prime = 18'b000000000010001001;
		14'b00111100011100:	sigmoid_prime = 18'b000000000010001001;
		14'b00111100011101:	sigmoid_prime = 18'b000000000010001000;
		14'b00111100011110:	sigmoid_prime = 18'b000000000010001000;
		14'b00111100011111:	sigmoid_prime = 18'b000000000010001000;
		14'b00111100100000:	sigmoid_prime = 18'b000000000010001000;
		14'b00111100100001:	sigmoid_prime = 18'b000000000010000111;
		14'b00111100100010:	sigmoid_prime = 18'b000000000010000111;
		14'b00111100100011:	sigmoid_prime = 18'b000000000010000111;
		14'b00111100100100:	sigmoid_prime = 18'b000000000010000111;
		14'b00111100100101:	sigmoid_prime = 18'b000000000010000110;
		14'b00111100100110:	sigmoid_prime = 18'b000000000010000110;
		14'b00111100100111:	sigmoid_prime = 18'b000000000010000110;
		14'b00111100101000:	sigmoid_prime = 18'b000000000010000101;
		14'b00111100101001:	sigmoid_prime = 18'b000000000010000101;
		14'b00111100101010:	sigmoid_prime = 18'b000000000010000101;
		14'b00111100101011:	sigmoid_prime = 18'b000000000010000101;
		14'b00111100101100:	sigmoid_prime = 18'b000000000010000100;
		14'b00111100101101:	sigmoid_prime = 18'b000000000010000100;
		14'b00111100101110:	sigmoid_prime = 18'b000000000010000100;
		14'b00111100101111:	sigmoid_prime = 18'b000000000010000100;
		14'b00111100110000:	sigmoid_prime = 18'b000000000010000011;
		14'b00111100110001:	sigmoid_prime = 18'b000000000010000011;
		14'b00111100110010:	sigmoid_prime = 18'b000000000010000011;
		14'b00111100110011:	sigmoid_prime = 18'b000000000010000011;
		14'b00111100110100:	sigmoid_prime = 18'b000000000010000010;
		14'b00111100110101:	sigmoid_prime = 18'b000000000010000010;
		14'b00111100110110:	sigmoid_prime = 18'b000000000010000010;
		14'b00111100110111:	sigmoid_prime = 18'b000000000010000010;
		14'b00111100111000:	sigmoid_prime = 18'b000000000010000001;
		14'b00111100111001:	sigmoid_prime = 18'b000000000010000001;
		14'b00111100111010:	sigmoid_prime = 18'b000000000010000001;
		14'b00111100111011:	sigmoid_prime = 18'b000000000010000001;
		14'b00111100111100:	sigmoid_prime = 18'b000000000010000000;
		14'b00111100111101:	sigmoid_prime = 18'b000000000010000000;
		14'b00111100111110:	sigmoid_prime = 18'b000000000010000000;
		14'b00111100111111:	sigmoid_prime = 18'b000000000010000000;
		14'b00111101000000:	sigmoid_prime = 18'b000000000001111111;
		14'b00111101000001:	sigmoid_prime = 18'b000000000001111111;
		14'b00111101000010:	sigmoid_prime = 18'b000000000001111111;
		14'b00111101000011:	sigmoid_prime = 18'b000000000001111111;
		14'b00111101000100:	sigmoid_prime = 18'b000000000001111110;
		14'b00111101000101:	sigmoid_prime = 18'b000000000001111110;
		14'b00111101000110:	sigmoid_prime = 18'b000000000001111110;
		14'b00111101000111:	sigmoid_prime = 18'b000000000001111110;
		14'b00111101001000:	sigmoid_prime = 18'b000000000001111101;
		14'b00111101001001:	sigmoid_prime = 18'b000000000001111101;
		14'b00111101001010:	sigmoid_prime = 18'b000000000001111101;
		14'b00111101001011:	sigmoid_prime = 18'b000000000001111101;
		14'b00111101001100:	sigmoid_prime = 18'b000000000001111100;
		14'b00111101001101:	sigmoid_prime = 18'b000000000001111100;
		14'b00111101001110:	sigmoid_prime = 18'b000000000001111100;
		14'b00111101001111:	sigmoid_prime = 18'b000000000001111100;
		14'b00111101010000:	sigmoid_prime = 18'b000000000001111011;
		14'b00111101010001:	sigmoid_prime = 18'b000000000001111011;
		14'b00111101010010:	sigmoid_prime = 18'b000000000001111011;
		14'b00111101010011:	sigmoid_prime = 18'b000000000001111011;
		14'b00111101010100:	sigmoid_prime = 18'b000000000001111010;
		14'b00111101010101:	sigmoid_prime = 18'b000000000001111010;
		14'b00111101010110:	sigmoid_prime = 18'b000000000001111010;
		14'b00111101010111:	sigmoid_prime = 18'b000000000001111010;
		14'b00111101011000:	sigmoid_prime = 18'b000000000001111001;
		14'b00111101011001:	sigmoid_prime = 18'b000000000001111001;
		14'b00111101011010:	sigmoid_prime = 18'b000000000001111001;
		14'b00111101011011:	sigmoid_prime = 18'b000000000001111001;
		14'b00111101011100:	sigmoid_prime = 18'b000000000001111001;
		14'b00111101011101:	sigmoid_prime = 18'b000000000001111000;
		14'b00111101011110:	sigmoid_prime = 18'b000000000001111000;
		14'b00111101011111:	sigmoid_prime = 18'b000000000001111000;
		14'b00111101100000:	sigmoid_prime = 18'b000000000001111000;
		14'b00111101100001:	sigmoid_prime = 18'b000000000001110111;
		14'b00111101100010:	sigmoid_prime = 18'b000000000001110111;
		14'b00111101100011:	sigmoid_prime = 18'b000000000001110111;
		14'b00111101100100:	sigmoid_prime = 18'b000000000001110111;
		14'b00111101100101:	sigmoid_prime = 18'b000000000001110110;
		14'b00111101100110:	sigmoid_prime = 18'b000000000001110110;
		14'b00111101100111:	sigmoid_prime = 18'b000000000001110110;
		14'b00111101101000:	sigmoid_prime = 18'b000000000001110110;
		14'b00111101101001:	sigmoid_prime = 18'b000000000001110101;
		14'b00111101101010:	sigmoid_prime = 18'b000000000001110101;
		14'b00111101101011:	sigmoid_prime = 18'b000000000001110101;
		14'b00111101101100:	sigmoid_prime = 18'b000000000001110101;
		14'b00111101101101:	sigmoid_prime = 18'b000000000001110101;
		14'b00111101101110:	sigmoid_prime = 18'b000000000001110100;
		14'b00111101101111:	sigmoid_prime = 18'b000000000001110100;
		14'b00111101110000:	sigmoid_prime = 18'b000000000001110100;
		14'b00111101110001:	sigmoid_prime = 18'b000000000001110100;
		14'b00111101110010:	sigmoid_prime = 18'b000000000001110011;
		14'b00111101110011:	sigmoid_prime = 18'b000000000001110011;
		14'b00111101110100:	sigmoid_prime = 18'b000000000001110011;
		14'b00111101110101:	sigmoid_prime = 18'b000000000001110011;
		14'b00111101110110:	sigmoid_prime = 18'b000000000001110011;
		14'b00111101110111:	sigmoid_prime = 18'b000000000001110010;
		14'b00111101111000:	sigmoid_prime = 18'b000000000001110010;
		14'b00111101111001:	sigmoid_prime = 18'b000000000001110010;
		14'b00111101111010:	sigmoid_prime = 18'b000000000001110010;
		14'b00111101111011:	sigmoid_prime = 18'b000000000001110001;
		14'b00111101111100:	sigmoid_prime = 18'b000000000001110001;
		14'b00111101111101:	sigmoid_prime = 18'b000000000001110001;
		14'b00111101111110:	sigmoid_prime = 18'b000000000001110001;
		14'b00111101111111:	sigmoid_prime = 18'b000000000001110001;
		14'b00111110000000:	sigmoid_prime = 18'b000000000001110000;
		14'b00111110000001:	sigmoid_prime = 18'b000000000001110000;
		14'b00111110000010:	sigmoid_prime = 18'b000000000001110000;
		14'b00111110000011:	sigmoid_prime = 18'b000000000001110000;
		14'b00111110000100:	sigmoid_prime = 18'b000000000001101111;
		14'b00111110000101:	sigmoid_prime = 18'b000000000001101111;
		14'b00111110000110:	sigmoid_prime = 18'b000000000001101111;
		14'b00111110000111:	sigmoid_prime = 18'b000000000001101111;
		14'b00111110001000:	sigmoid_prime = 18'b000000000001101111;
		14'b00111110001001:	sigmoid_prime = 18'b000000000001101110;
		14'b00111110001010:	sigmoid_prime = 18'b000000000001101110;
		14'b00111110001011:	sigmoid_prime = 18'b000000000001101110;
		14'b00111110001100:	sigmoid_prime = 18'b000000000001101110;
		14'b00111110001101:	sigmoid_prime = 18'b000000000001101101;
		14'b00111110001110:	sigmoid_prime = 18'b000000000001101101;
		14'b00111110001111:	sigmoid_prime = 18'b000000000001101101;
		14'b00111110010000:	sigmoid_prime = 18'b000000000001101101;
		14'b00111110010001:	sigmoid_prime = 18'b000000000001101101;
		14'b00111110010010:	sigmoid_prime = 18'b000000000001101100;
		14'b00111110010011:	sigmoid_prime = 18'b000000000001101100;
		14'b00111110010100:	sigmoid_prime = 18'b000000000001101100;
		14'b00111110010101:	sigmoid_prime = 18'b000000000001101100;
		14'b00111110010110:	sigmoid_prime = 18'b000000000001101100;
		14'b00111110010111:	sigmoid_prime = 18'b000000000001101011;
		14'b00111110011000:	sigmoid_prime = 18'b000000000001101011;
		14'b00111110011001:	sigmoid_prime = 18'b000000000001101011;
		14'b00111110011010:	sigmoid_prime = 18'b000000000001101011;
		14'b00111110011011:	sigmoid_prime = 18'b000000000001101011;
		14'b00111110011100:	sigmoid_prime = 18'b000000000001101010;
		14'b00111110011101:	sigmoid_prime = 18'b000000000001101010;
		14'b00111110011110:	sigmoid_prime = 18'b000000000001101010;
		14'b00111110011111:	sigmoid_prime = 18'b000000000001101010;
		14'b00111110100000:	sigmoid_prime = 18'b000000000001101001;
		14'b00111110100001:	sigmoid_prime = 18'b000000000001101001;
		14'b00111110100010:	sigmoid_prime = 18'b000000000001101001;
		14'b00111110100011:	sigmoid_prime = 18'b000000000001101001;
		14'b00111110100100:	sigmoid_prime = 18'b000000000001101001;
		14'b00111110100101:	sigmoid_prime = 18'b000000000001101000;
		14'b00111110100110:	sigmoid_prime = 18'b000000000001101000;
		14'b00111110100111:	sigmoid_prime = 18'b000000000001101000;
		14'b00111110101000:	sigmoid_prime = 18'b000000000001101000;
		14'b00111110101001:	sigmoid_prime = 18'b000000000001101000;
		14'b00111110101010:	sigmoid_prime = 18'b000000000001100111;
		14'b00111110101011:	sigmoid_prime = 18'b000000000001100111;
		14'b00111110101100:	sigmoid_prime = 18'b000000000001100111;
		14'b00111110101101:	sigmoid_prime = 18'b000000000001100111;
		14'b00111110101110:	sigmoid_prime = 18'b000000000001100111;
		14'b00111110101111:	sigmoid_prime = 18'b000000000001100110;
		14'b00111110110000:	sigmoid_prime = 18'b000000000001100110;
		14'b00111110110001:	sigmoid_prime = 18'b000000000001100110;
		14'b00111110110010:	sigmoid_prime = 18'b000000000001100110;
		14'b00111110110011:	sigmoid_prime = 18'b000000000001100110;
		14'b00111110110100:	sigmoid_prime = 18'b000000000001100101;
		14'b00111110110101:	sigmoid_prime = 18'b000000000001100101;
		14'b00111110110110:	sigmoid_prime = 18'b000000000001100101;
		14'b00111110110111:	sigmoid_prime = 18'b000000000001100101;
		14'b00111110111000:	sigmoid_prime = 18'b000000000001100101;
		14'b00111110111001:	sigmoid_prime = 18'b000000000001100100;
		14'b00111110111010:	sigmoid_prime = 18'b000000000001100100;
		14'b00111110111011:	sigmoid_prime = 18'b000000000001100100;
		14'b00111110111100:	sigmoid_prime = 18'b000000000001100100;
		14'b00111110111101:	sigmoid_prime = 18'b000000000001100100;
		14'b00111110111110:	sigmoid_prime = 18'b000000000001100011;
		14'b00111110111111:	sigmoid_prime = 18'b000000000001100011;
		14'b00111111000000:	sigmoid_prime = 18'b000000000001100011;
		14'b00111111000001:	sigmoid_prime = 18'b000000000001100011;
		14'b00111111000010:	sigmoid_prime = 18'b000000000001100011;
		14'b00111111000011:	sigmoid_prime = 18'b000000000001100010;
		14'b00111111000100:	sigmoid_prime = 18'b000000000001100010;
		14'b00111111000101:	sigmoid_prime = 18'b000000000001100010;
		14'b00111111000110:	sigmoid_prime = 18'b000000000001100010;
		14'b00111111000111:	sigmoid_prime = 18'b000000000001100010;
		14'b00111111001000:	sigmoid_prime = 18'b000000000001100010;
		14'b00111111001001:	sigmoid_prime = 18'b000000000001100001;
		14'b00111111001010:	sigmoid_prime = 18'b000000000001100001;
		14'b00111111001011:	sigmoid_prime = 18'b000000000001100001;
		14'b00111111001100:	sigmoid_prime = 18'b000000000001100001;
		14'b00111111001101:	sigmoid_prime = 18'b000000000001100001;
		14'b00111111001110:	sigmoid_prime = 18'b000000000001100000;
		14'b00111111001111:	sigmoid_prime = 18'b000000000001100000;
		14'b00111111010000:	sigmoid_prime = 18'b000000000001100000;
		14'b00111111010001:	sigmoid_prime = 18'b000000000001100000;
		14'b00111111010010:	sigmoid_prime = 18'b000000000001100000;
		14'b00111111010011:	sigmoid_prime = 18'b000000000001011111;
		14'b00111111010100:	sigmoid_prime = 18'b000000000001011111;
		14'b00111111010101:	sigmoid_prime = 18'b000000000001011111;
		14'b00111111010110:	sigmoid_prime = 18'b000000000001011111;
		14'b00111111010111:	sigmoid_prime = 18'b000000000001011111;
		14'b00111111011000:	sigmoid_prime = 18'b000000000001011111;
		14'b00111111011001:	sigmoid_prime = 18'b000000000001011110;
		14'b00111111011010:	sigmoid_prime = 18'b000000000001011110;
		14'b00111111011011:	sigmoid_prime = 18'b000000000001011110;
		14'b00111111011100:	sigmoid_prime = 18'b000000000001011110;
		14'b00111111011101:	sigmoid_prime = 18'b000000000001011110;
		14'b00111111011110:	sigmoid_prime = 18'b000000000001011101;
		14'b00111111011111:	sigmoid_prime = 18'b000000000001011101;
		14'b00111111100000:	sigmoid_prime = 18'b000000000001011101;
		14'b00111111100001:	sigmoid_prime = 18'b000000000001011101;
		14'b00111111100010:	sigmoid_prime = 18'b000000000001011101;
		14'b00111111100011:	sigmoid_prime = 18'b000000000001011100;
		14'b00111111100100:	sigmoid_prime = 18'b000000000001011100;
		14'b00111111100101:	sigmoid_prime = 18'b000000000001011100;
		14'b00111111100110:	sigmoid_prime = 18'b000000000001011100;
		14'b00111111100111:	sigmoid_prime = 18'b000000000001011100;
		14'b00111111101000:	sigmoid_prime = 18'b000000000001011100;
		14'b00111111101001:	sigmoid_prime = 18'b000000000001011011;
		14'b00111111101010:	sigmoid_prime = 18'b000000000001011011;
		14'b00111111101011:	sigmoid_prime = 18'b000000000001011011;
		14'b00111111101100:	sigmoid_prime = 18'b000000000001011011;
		14'b00111111101101:	sigmoid_prime = 18'b000000000001011011;
		14'b00111111101110:	sigmoid_prime = 18'b000000000001011011;
		14'b00111111101111:	sigmoid_prime = 18'b000000000001011010;
		14'b00111111110000:	sigmoid_prime = 18'b000000000001011010;
		14'b00111111110001:	sigmoid_prime = 18'b000000000001011010;
		14'b00111111110010:	sigmoid_prime = 18'b000000000001011010;
		14'b00111111110011:	sigmoid_prime = 18'b000000000001011010;
		14'b00111111110100:	sigmoid_prime = 18'b000000000001011001;
		14'b00111111110101:	sigmoid_prime = 18'b000000000001011001;
		14'b00111111110110:	sigmoid_prime = 18'b000000000001011001;
		14'b00111111110111:	sigmoid_prime = 18'b000000000001011001;
		14'b00111111111000:	sigmoid_prime = 18'b000000000001011001;
		14'b00111111111001:	sigmoid_prime = 18'b000000000001011001;
		14'b00111111111010:	sigmoid_prime = 18'b000000000001011000;
		14'b00111111111011:	sigmoid_prime = 18'b000000000001011000;
		14'b00111111111100:	sigmoid_prime = 18'b000000000001011000;
		14'b00111111111101:	sigmoid_prime = 18'b000000000001011000;
		14'b00111111111110:	sigmoid_prime = 18'b000000000001011000;
		14'b00111111111111:	sigmoid_prime = 18'b000000000001011000;
		14'b01000000000000:	sigmoid_prime = 18'b000000000001010111;
		14'b01000000000001:	sigmoid_prime = 18'b000000000001010111;
		14'b01000000000010:	sigmoid_prime = 18'b000000000001010111;
		14'b01000000000011:	sigmoid_prime = 18'b000000000001010111;
		14'b01000000000100:	sigmoid_prime = 18'b000000000001010111;
		14'b01000000000101:	sigmoid_prime = 18'b000000000001010111;
		14'b01000000000110:	sigmoid_prime = 18'b000000000001010110;
		14'b01000000000111:	sigmoid_prime = 18'b000000000001010110;
		14'b01000000001000:	sigmoid_prime = 18'b000000000001010110;
		14'b01000000001001:	sigmoid_prime = 18'b000000000001010110;
		14'b01000000001010:	sigmoid_prime = 18'b000000000001010110;
		14'b01000000001011:	sigmoid_prime = 18'b000000000001010110;
		14'b01000000001100:	sigmoid_prime = 18'b000000000001010101;
		14'b01000000001101:	sigmoid_prime = 18'b000000000001010101;
		14'b01000000001110:	sigmoid_prime = 18'b000000000001010101;
		14'b01000000001111:	sigmoid_prime = 18'b000000000001010101;
		14'b01000000010000:	sigmoid_prime = 18'b000000000001010101;
		14'b01000000010001:	sigmoid_prime = 18'b000000000001010101;
		14'b01000000010010:	sigmoid_prime = 18'b000000000001010100;
		14'b01000000010011:	sigmoid_prime = 18'b000000000001010100;
		14'b01000000010100:	sigmoid_prime = 18'b000000000001010100;
		14'b01000000010101:	sigmoid_prime = 18'b000000000001010100;
		14'b01000000010110:	sigmoid_prime = 18'b000000000001010100;
		14'b01000000010111:	sigmoid_prime = 18'b000000000001010100;
		14'b01000000011000:	sigmoid_prime = 18'b000000000001010011;
		14'b01000000011001:	sigmoid_prime = 18'b000000000001010011;
		14'b01000000011010:	sigmoid_prime = 18'b000000000001010011;
		14'b01000000011011:	sigmoid_prime = 18'b000000000001010011;
		14'b01000000011100:	sigmoid_prime = 18'b000000000001010011;
		14'b01000000011101:	sigmoid_prime = 18'b000000000001010011;
		14'b01000000011110:	sigmoid_prime = 18'b000000000001010010;
		14'b01000000011111:	sigmoid_prime = 18'b000000000001010010;
		14'b01000000100000:	sigmoid_prime = 18'b000000000001010010;
		14'b01000000100001:	sigmoid_prime = 18'b000000000001010010;
		14'b01000000100010:	sigmoid_prime = 18'b000000000001010010;
		14'b01000000100011:	sigmoid_prime = 18'b000000000001010010;
		14'b01000000100100:	sigmoid_prime = 18'b000000000001010001;
		14'b01000000100101:	sigmoid_prime = 18'b000000000001010001;
		14'b01000000100110:	sigmoid_prime = 18'b000000000001010001;
		14'b01000000100111:	sigmoid_prime = 18'b000000000001010001;
		14'b01000000101000:	sigmoid_prime = 18'b000000000001010001;
		14'b01000000101001:	sigmoid_prime = 18'b000000000001010001;
		14'b01000000101010:	sigmoid_prime = 18'b000000000001010000;
		14'b01000000101011:	sigmoid_prime = 18'b000000000001010000;
		14'b01000000101100:	sigmoid_prime = 18'b000000000001010000;
		14'b01000000101101:	sigmoid_prime = 18'b000000000001010000;
		14'b01000000101110:	sigmoid_prime = 18'b000000000001010000;
		14'b01000000101111:	sigmoid_prime = 18'b000000000001010000;
		14'b01000000110000:	sigmoid_prime = 18'b000000000001010000;
		14'b01000000110001:	sigmoid_prime = 18'b000000000001001111;
		14'b01000000110010:	sigmoid_prime = 18'b000000000001001111;
		14'b01000000110011:	sigmoid_prime = 18'b000000000001001111;
		14'b01000000110100:	sigmoid_prime = 18'b000000000001001111;
		14'b01000000110101:	sigmoid_prime = 18'b000000000001001111;
		14'b01000000110110:	sigmoid_prime = 18'b000000000001001111;
		14'b01000000110111:	sigmoid_prime = 18'b000000000001001110;
		14'b01000000111000:	sigmoid_prime = 18'b000000000001001110;
		14'b01000000111001:	sigmoid_prime = 18'b000000000001001110;
		14'b01000000111010:	sigmoid_prime = 18'b000000000001001110;
		14'b01000000111011:	sigmoid_prime = 18'b000000000001001110;
		14'b01000000111100:	sigmoid_prime = 18'b000000000001001110;
		14'b01000000111101:	sigmoid_prime = 18'b000000000001001110;
		14'b01000000111110:	sigmoid_prime = 18'b000000000001001101;
		14'b01000000111111:	sigmoid_prime = 18'b000000000001001101;
		14'b01000001000000:	sigmoid_prime = 18'b000000000001001101;
		14'b01000001000001:	sigmoid_prime = 18'b000000000001001101;
		14'b01000001000010:	sigmoid_prime = 18'b000000000001001101;
		14'b01000001000011:	sigmoid_prime = 18'b000000000001001101;
		14'b01000001000100:	sigmoid_prime = 18'b000000000001001100;
		14'b01000001000101:	sigmoid_prime = 18'b000000000001001100;
		14'b01000001000110:	sigmoid_prime = 18'b000000000001001100;
		14'b01000001000111:	sigmoid_prime = 18'b000000000001001100;
		14'b01000001001000:	sigmoid_prime = 18'b000000000001001100;
		14'b01000001001001:	sigmoid_prime = 18'b000000000001001100;
		14'b01000001001010:	sigmoid_prime = 18'b000000000001001100;
		14'b01000001001011:	sigmoid_prime = 18'b000000000001001011;
		14'b01000001001100:	sigmoid_prime = 18'b000000000001001011;
		14'b01000001001101:	sigmoid_prime = 18'b000000000001001011;
		14'b01000001001110:	sigmoid_prime = 18'b000000000001001011;
		14'b01000001001111:	sigmoid_prime = 18'b000000000001001011;
		14'b01000001010000:	sigmoid_prime = 18'b000000000001001011;
		14'b01000001010001:	sigmoid_prime = 18'b000000000001001011;
		14'b01000001010010:	sigmoid_prime = 18'b000000000001001010;
		14'b01000001010011:	sigmoid_prime = 18'b000000000001001010;
		14'b01000001010100:	sigmoid_prime = 18'b000000000001001010;
		14'b01000001010101:	sigmoid_prime = 18'b000000000001001010;
		14'b01000001010110:	sigmoid_prime = 18'b000000000001001010;
		14'b01000001010111:	sigmoid_prime = 18'b000000000001001010;
		14'b01000001011000:	sigmoid_prime = 18'b000000000001001010;
		14'b01000001011001:	sigmoid_prime = 18'b000000000001001001;
		14'b01000001011010:	sigmoid_prime = 18'b000000000001001001;
		14'b01000001011011:	sigmoid_prime = 18'b000000000001001001;
		14'b01000001011100:	sigmoid_prime = 18'b000000000001001001;
		14'b01000001011101:	sigmoid_prime = 18'b000000000001001001;
		14'b01000001011110:	sigmoid_prime = 18'b000000000001001001;
		14'b01000001011111:	sigmoid_prime = 18'b000000000001001001;
		14'b01000001100000:	sigmoid_prime = 18'b000000000001001000;
		14'b01000001100001:	sigmoid_prime = 18'b000000000001001000;
		14'b01000001100010:	sigmoid_prime = 18'b000000000001001000;
		14'b01000001100011:	sigmoid_prime = 18'b000000000001001000;
		14'b01000001100100:	sigmoid_prime = 18'b000000000001001000;
		14'b01000001100101:	sigmoid_prime = 18'b000000000001001000;
		14'b01000001100110:	sigmoid_prime = 18'b000000000001001000;
		14'b01000001100111:	sigmoid_prime = 18'b000000000001000111;
		14'b01000001101000:	sigmoid_prime = 18'b000000000001000111;
		14'b01000001101001:	sigmoid_prime = 18'b000000000001000111;
		14'b01000001101010:	sigmoid_prime = 18'b000000000001000111;
		14'b01000001101011:	sigmoid_prime = 18'b000000000001000111;
		14'b01000001101100:	sigmoid_prime = 18'b000000000001000111;
		14'b01000001101101:	sigmoid_prime = 18'b000000000001000111;
		14'b01000001101110:	sigmoid_prime = 18'b000000000001000110;
		14'b01000001101111:	sigmoid_prime = 18'b000000000001000110;
		14'b01000001110000:	sigmoid_prime = 18'b000000000001000110;
		14'b01000001110001:	sigmoid_prime = 18'b000000000001000110;
		14'b01000001110010:	sigmoid_prime = 18'b000000000001000110;
		14'b01000001110011:	sigmoid_prime = 18'b000000000001000110;
		14'b01000001110100:	sigmoid_prime = 18'b000000000001000110;
		14'b01000001110101:	sigmoid_prime = 18'b000000000001000101;
		14'b01000001110110:	sigmoid_prime = 18'b000000000001000101;
		14'b01000001110111:	sigmoid_prime = 18'b000000000001000101;
		14'b01000001111000:	sigmoid_prime = 18'b000000000001000101;
		14'b01000001111001:	sigmoid_prime = 18'b000000000001000101;
		14'b01000001111010:	sigmoid_prime = 18'b000000000001000101;
		14'b01000001111011:	sigmoid_prime = 18'b000000000001000101;
		14'b01000001111100:	sigmoid_prime = 18'b000000000001000100;
		14'b01000001111101:	sigmoid_prime = 18'b000000000001000100;
		14'b01000001111110:	sigmoid_prime = 18'b000000000001000100;
		14'b01000001111111:	sigmoid_prime = 18'b000000000001000100;
		14'b01000010000000:	sigmoid_prime = 18'b000000000001000100;
		14'b01000010000001:	sigmoid_prime = 18'b000000000001000100;
		14'b01000010000010:	sigmoid_prime = 18'b000000000001000100;
		14'b01000010000011:	sigmoid_prime = 18'b000000000001000100;
		14'b01000010000100:	sigmoid_prime = 18'b000000000001000011;
		14'b01000010000101:	sigmoid_prime = 18'b000000000001000011;
		14'b01000010000110:	sigmoid_prime = 18'b000000000001000011;
		14'b01000010000111:	sigmoid_prime = 18'b000000000001000011;
		14'b01000010001000:	sigmoid_prime = 18'b000000000001000011;
		14'b01000010001001:	sigmoid_prime = 18'b000000000001000011;
		14'b01000010001010:	sigmoid_prime = 18'b000000000001000011;
		14'b01000010001011:	sigmoid_prime = 18'b000000000001000010;
		14'b01000010001100:	sigmoid_prime = 18'b000000000001000010;
		14'b01000010001101:	sigmoid_prime = 18'b000000000001000010;
		14'b01000010001110:	sigmoid_prime = 18'b000000000001000010;
		14'b01000010001111:	sigmoid_prime = 18'b000000000001000010;
		14'b01000010010000:	sigmoid_prime = 18'b000000000001000010;
		14'b01000010010001:	sigmoid_prime = 18'b000000000001000010;
		14'b01000010010010:	sigmoid_prime = 18'b000000000001000010;
		14'b01000010010011:	sigmoid_prime = 18'b000000000001000001;
		14'b01000010010100:	sigmoid_prime = 18'b000000000001000001;
		14'b01000010010101:	sigmoid_prime = 18'b000000000001000001;
		14'b01000010010110:	sigmoid_prime = 18'b000000000001000001;
		14'b01000010010111:	sigmoid_prime = 18'b000000000001000001;
		14'b01000010011000:	sigmoid_prime = 18'b000000000001000001;
		14'b01000010011001:	sigmoid_prime = 18'b000000000001000001;
		14'b01000010011010:	sigmoid_prime = 18'b000000000001000001;
		14'b01000010011011:	sigmoid_prime = 18'b000000000001000000;
		14'b01000010011100:	sigmoid_prime = 18'b000000000001000000;
		14'b01000010011101:	sigmoid_prime = 18'b000000000001000000;
		14'b01000010011110:	sigmoid_prime = 18'b000000000001000000;
		14'b01000010011111:	sigmoid_prime = 18'b000000000001000000;
		14'b01000010100000:	sigmoid_prime = 18'b000000000001000000;
		14'b01000010100001:	sigmoid_prime = 18'b000000000001000000;
		14'b01000010100010:	sigmoid_prime = 18'b000000000001000000;
		14'b01000010100011:	sigmoid_prime = 18'b000000000000111111;
		14'b01000010100100:	sigmoid_prime = 18'b000000000000111111;
		14'b01000010100101:	sigmoid_prime = 18'b000000000000111111;
		14'b01000010100110:	sigmoid_prime = 18'b000000000000111111;
		14'b01000010100111:	sigmoid_prime = 18'b000000000000111111;
		14'b01000010101000:	sigmoid_prime = 18'b000000000000111111;
		14'b01000010101001:	sigmoid_prime = 18'b000000000000111111;
		14'b01000010101010:	sigmoid_prime = 18'b000000000000111111;
		14'b01000010101011:	sigmoid_prime = 18'b000000000000111110;
		14'b01000010101100:	sigmoid_prime = 18'b000000000000111110;
		14'b01000010101101:	sigmoid_prime = 18'b000000000000111110;
		14'b01000010101110:	sigmoid_prime = 18'b000000000000111110;
		14'b01000010101111:	sigmoid_prime = 18'b000000000000111110;
		14'b01000010110000:	sigmoid_prime = 18'b000000000000111110;
		14'b01000010110001:	sigmoid_prime = 18'b000000000000111110;
		14'b01000010110010:	sigmoid_prime = 18'b000000000000111110;
		14'b01000010110011:	sigmoid_prime = 18'b000000000000111101;
		14'b01000010110100:	sigmoid_prime = 18'b000000000000111101;
		14'b01000010110101:	sigmoid_prime = 18'b000000000000111101;
		14'b01000010110110:	sigmoid_prime = 18'b000000000000111101;
		14'b01000010110111:	sigmoid_prime = 18'b000000000000111101;
		14'b01000010111000:	sigmoid_prime = 18'b000000000000111101;
		14'b01000010111001:	sigmoid_prime = 18'b000000000000111101;
		14'b01000010111010:	sigmoid_prime = 18'b000000000000111101;
		14'b01000010111011:	sigmoid_prime = 18'b000000000000111101;
		14'b01000010111100:	sigmoid_prime = 18'b000000000000111100;
		14'b01000010111101:	sigmoid_prime = 18'b000000000000111100;
		14'b01000010111110:	sigmoid_prime = 18'b000000000000111100;
		14'b01000010111111:	sigmoid_prime = 18'b000000000000111100;
		14'b01000011000000:	sigmoid_prime = 18'b000000000000111100;
		14'b01000011000001:	sigmoid_prime = 18'b000000000000111100;
		14'b01000011000010:	sigmoid_prime = 18'b000000000000111100;
		14'b01000011000011:	sigmoid_prime = 18'b000000000000111100;
		14'b01000011000100:	sigmoid_prime = 18'b000000000000111011;
		14'b01000011000101:	sigmoid_prime = 18'b000000000000111011;
		14'b01000011000110:	sigmoid_prime = 18'b000000000000111011;
		14'b01000011000111:	sigmoid_prime = 18'b000000000000111011;
		14'b01000011001000:	sigmoid_prime = 18'b000000000000111011;
		14'b01000011001001:	sigmoid_prime = 18'b000000000000111011;
		14'b01000011001010:	sigmoid_prime = 18'b000000000000111011;
		14'b01000011001011:	sigmoid_prime = 18'b000000000000111011;
		14'b01000011001100:	sigmoid_prime = 18'b000000000000111011;
		14'b01000011001101:	sigmoid_prime = 18'b000000000000111010;
		14'b01000011001110:	sigmoid_prime = 18'b000000000000111010;
		14'b01000011001111:	sigmoid_prime = 18'b000000000000111010;
		14'b01000011010000:	sigmoid_prime = 18'b000000000000111010;
		14'b01000011010001:	sigmoid_prime = 18'b000000000000111010;
		14'b01000011010010:	sigmoid_prime = 18'b000000000000111010;
		14'b01000011010011:	sigmoid_prime = 18'b000000000000111010;
		14'b01000011010100:	sigmoid_prime = 18'b000000000000111010;
		14'b01000011010101:	sigmoid_prime = 18'b000000000000111001;
		14'b01000011010110:	sigmoid_prime = 18'b000000000000111001;
		14'b01000011010111:	sigmoid_prime = 18'b000000000000111001;
		14'b01000011011000:	sigmoid_prime = 18'b000000000000111001;
		14'b01000011011001:	sigmoid_prime = 18'b000000000000111001;
		14'b01000011011010:	sigmoid_prime = 18'b000000000000111001;
		14'b01000011011011:	sigmoid_prime = 18'b000000000000111001;
		14'b01000011011100:	sigmoid_prime = 18'b000000000000111001;
		14'b01000011011101:	sigmoid_prime = 18'b000000000000111001;
		14'b01000011011110:	sigmoid_prime = 18'b000000000000111000;
		14'b01000011011111:	sigmoid_prime = 18'b000000000000111000;
		14'b01000011100000:	sigmoid_prime = 18'b000000000000111000;
		14'b01000011100001:	sigmoid_prime = 18'b000000000000111000;
		14'b01000011100010:	sigmoid_prime = 18'b000000000000111000;
		14'b01000011100011:	sigmoid_prime = 18'b000000000000111000;
		14'b01000011100100:	sigmoid_prime = 18'b000000000000111000;
		14'b01000011100101:	sigmoid_prime = 18'b000000000000111000;
		14'b01000011100110:	sigmoid_prime = 18'b000000000000111000;
		14'b01000011100111:	sigmoid_prime = 18'b000000000000110111;
		14'b01000011101000:	sigmoid_prime = 18'b000000000000110111;
		14'b01000011101001:	sigmoid_prime = 18'b000000000000110111;
		14'b01000011101010:	sigmoid_prime = 18'b000000000000110111;
		14'b01000011101011:	sigmoid_prime = 18'b000000000000110111;
		14'b01000011101100:	sigmoid_prime = 18'b000000000000110111;
		14'b01000011101101:	sigmoid_prime = 18'b000000000000110111;
		14'b01000011101110:	sigmoid_prime = 18'b000000000000110111;
		14'b01000011101111:	sigmoid_prime = 18'b000000000000110111;
		14'b01000011110000:	sigmoid_prime = 18'b000000000000110111;
		14'b01000011110001:	sigmoid_prime = 18'b000000000000110110;
		14'b01000011110010:	sigmoid_prime = 18'b000000000000110110;
		14'b01000011110011:	sigmoid_prime = 18'b000000000000110110;
		14'b01000011110100:	sigmoid_prime = 18'b000000000000110110;
		14'b01000011110101:	sigmoid_prime = 18'b000000000000110110;
		14'b01000011110110:	sigmoid_prime = 18'b000000000000110110;
		14'b01000011110111:	sigmoid_prime = 18'b000000000000110110;
		14'b01000011111000:	sigmoid_prime = 18'b000000000000110110;
		14'b01000011111001:	sigmoid_prime = 18'b000000000000110110;
		14'b01000011111010:	sigmoid_prime = 18'b000000000000110101;
		14'b01000011111011:	sigmoid_prime = 18'b000000000000110101;
		14'b01000011111100:	sigmoid_prime = 18'b000000000000110101;
		14'b01000011111101:	sigmoid_prime = 18'b000000000000110101;
		14'b01000011111110:	sigmoid_prime = 18'b000000000000110101;
		14'b01000011111111:	sigmoid_prime = 18'b000000000000110101;
		14'b01000100000000:	sigmoid_prime = 18'b000000000000110101;
		14'b01000100000001:	sigmoid_prime = 18'b000000000000110101;
		14'b01000100000010:	sigmoid_prime = 18'b000000000000110101;
		14'b01000100000011:	sigmoid_prime = 18'b000000000000110101;
		14'b01000100000100:	sigmoid_prime = 18'b000000000000110100;
		14'b01000100000101:	sigmoid_prime = 18'b000000000000110100;
		14'b01000100000110:	sigmoid_prime = 18'b000000000000110100;
		14'b01000100000111:	sigmoid_prime = 18'b000000000000110100;
		14'b01000100001000:	sigmoid_prime = 18'b000000000000110100;
		14'b01000100001001:	sigmoid_prime = 18'b000000000000110100;
		14'b01000100001010:	sigmoid_prime = 18'b000000000000110100;
		14'b01000100001011:	sigmoid_prime = 18'b000000000000110100;
		14'b01000100001100:	sigmoid_prime = 18'b000000000000110100;
		14'b01000100001101:	sigmoid_prime = 18'b000000000000110011;
		14'b01000100001110:	sigmoid_prime = 18'b000000000000110011;
		14'b01000100001111:	sigmoid_prime = 18'b000000000000110011;
		14'b01000100010000:	sigmoid_prime = 18'b000000000000110011;
		14'b01000100010001:	sigmoid_prime = 18'b000000000000110011;
		14'b01000100010010:	sigmoid_prime = 18'b000000000000110011;
		14'b01000100010011:	sigmoid_prime = 18'b000000000000110011;
		14'b01000100010100:	sigmoid_prime = 18'b000000000000110011;
		14'b01000100010101:	sigmoid_prime = 18'b000000000000110011;
		14'b01000100010110:	sigmoid_prime = 18'b000000000000110011;
		14'b01000100010111:	sigmoid_prime = 18'b000000000000110010;
		14'b01000100011000:	sigmoid_prime = 18'b000000000000110010;
		14'b01000100011001:	sigmoid_prime = 18'b000000000000110010;
		14'b01000100011010:	sigmoid_prime = 18'b000000000000110010;
		14'b01000100011011:	sigmoid_prime = 18'b000000000000110010;
		14'b01000100011100:	sigmoid_prime = 18'b000000000000110010;
		14'b01000100011101:	sigmoid_prime = 18'b000000000000110010;
		14'b01000100011110:	sigmoid_prime = 18'b000000000000110010;
		14'b01000100011111:	sigmoid_prime = 18'b000000000000110010;
		14'b01000100100000:	sigmoid_prime = 18'b000000000000110010;
		14'b01000100100001:	sigmoid_prime = 18'b000000000000110001;
		14'b01000100100010:	sigmoid_prime = 18'b000000000000110001;
		14'b01000100100011:	sigmoid_prime = 18'b000000000000110001;
		14'b01000100100100:	sigmoid_prime = 18'b000000000000110001;
		14'b01000100100101:	sigmoid_prime = 18'b000000000000110001;
		14'b01000100100110:	sigmoid_prime = 18'b000000000000110001;
		14'b01000100100111:	sigmoid_prime = 18'b000000000000110001;
		14'b01000100101000:	sigmoid_prime = 18'b000000000000110001;
		14'b01000100101001:	sigmoid_prime = 18'b000000000000110001;
		14'b01000100101010:	sigmoid_prime = 18'b000000000000110001;
		14'b01000100101011:	sigmoid_prime = 18'b000000000000110001;
		14'b01000100101100:	sigmoid_prime = 18'b000000000000110000;
		14'b01000100101101:	sigmoid_prime = 18'b000000000000110000;
		14'b01000100101110:	sigmoid_prime = 18'b000000000000110000;
		14'b01000100101111:	sigmoid_prime = 18'b000000000000110000;
		14'b01000100110000:	sigmoid_prime = 18'b000000000000110000;
		14'b01000100110001:	sigmoid_prime = 18'b000000000000110000;
		14'b01000100110010:	sigmoid_prime = 18'b000000000000110000;
		14'b01000100110011:	sigmoid_prime = 18'b000000000000110000;
		14'b01000100110100:	sigmoid_prime = 18'b000000000000110000;
		14'b01000100110101:	sigmoid_prime = 18'b000000000000110000;
		14'b01000100110110:	sigmoid_prime = 18'b000000000000101111;
		14'b01000100110111:	sigmoid_prime = 18'b000000000000101111;
		14'b01000100111000:	sigmoid_prime = 18'b000000000000101111;
		14'b01000100111001:	sigmoid_prime = 18'b000000000000101111;
		14'b01000100111010:	sigmoid_prime = 18'b000000000000101111;
		14'b01000100111011:	sigmoid_prime = 18'b000000000000101111;
		14'b01000100111100:	sigmoid_prime = 18'b000000000000101111;
		14'b01000100111101:	sigmoid_prime = 18'b000000000000101111;
		14'b01000100111110:	sigmoid_prime = 18'b000000000000101111;
		14'b01000100111111:	sigmoid_prime = 18'b000000000000101111;
		14'b01000101000000:	sigmoid_prime = 18'b000000000000101111;
		14'b01000101000001:	sigmoid_prime = 18'b000000000000101110;
		14'b01000101000010:	sigmoid_prime = 18'b000000000000101110;
		14'b01000101000011:	sigmoid_prime = 18'b000000000000101110;
		14'b01000101000100:	sigmoid_prime = 18'b000000000000101110;
		14'b01000101000101:	sigmoid_prime = 18'b000000000000101110;
		14'b01000101000110:	sigmoid_prime = 18'b000000000000101110;
		14'b01000101000111:	sigmoid_prime = 18'b000000000000101110;
		14'b01000101001000:	sigmoid_prime = 18'b000000000000101110;
		14'b01000101001001:	sigmoid_prime = 18'b000000000000101110;
		14'b01000101001010:	sigmoid_prime = 18'b000000000000101110;
		14'b01000101001011:	sigmoid_prime = 18'b000000000000101110;
		14'b01000101001100:	sigmoid_prime = 18'b000000000000101101;
		14'b01000101001101:	sigmoid_prime = 18'b000000000000101101;
		14'b01000101001110:	sigmoid_prime = 18'b000000000000101101;
		14'b01000101001111:	sigmoid_prime = 18'b000000000000101101;
		14'b01000101010000:	sigmoid_prime = 18'b000000000000101101;
		14'b01000101010001:	sigmoid_prime = 18'b000000000000101101;
		14'b01000101010010:	sigmoid_prime = 18'b000000000000101101;
		14'b01000101010011:	sigmoid_prime = 18'b000000000000101101;
		14'b01000101010100:	sigmoid_prime = 18'b000000000000101101;
		14'b01000101010101:	sigmoid_prime = 18'b000000000000101101;
		14'b01000101010110:	sigmoid_prime = 18'b000000000000101101;
		14'b01000101010111:	sigmoid_prime = 18'b000000000000101100;
		14'b01000101011000:	sigmoid_prime = 18'b000000000000101100;
		14'b01000101011001:	sigmoid_prime = 18'b000000000000101100;
		14'b01000101011010:	sigmoid_prime = 18'b000000000000101100;
		14'b01000101011011:	sigmoid_prime = 18'b000000000000101100;
		14'b01000101011100:	sigmoid_prime = 18'b000000000000101100;
		14'b01000101011101:	sigmoid_prime = 18'b000000000000101100;
		14'b01000101011110:	sigmoid_prime = 18'b000000000000101100;
		14'b01000101011111:	sigmoid_prime = 18'b000000000000101100;
		14'b01000101100000:	sigmoid_prime = 18'b000000000000101100;
		14'b01000101100001:	sigmoid_prime = 18'b000000000000101100;
		14'b01000101100010:	sigmoid_prime = 18'b000000000000101100;
		14'b01000101100011:	sigmoid_prime = 18'b000000000000101011;
		14'b01000101100100:	sigmoid_prime = 18'b000000000000101011;
		14'b01000101100101:	sigmoid_prime = 18'b000000000000101011;
		14'b01000101100110:	sigmoid_prime = 18'b000000000000101011;
		14'b01000101100111:	sigmoid_prime = 18'b000000000000101011;
		14'b01000101101000:	sigmoid_prime = 18'b000000000000101011;
		14'b01000101101001:	sigmoid_prime = 18'b000000000000101011;
		14'b01000101101010:	sigmoid_prime = 18'b000000000000101011;
		14'b01000101101011:	sigmoid_prime = 18'b000000000000101011;
		14'b01000101101100:	sigmoid_prime = 18'b000000000000101011;
		14'b01000101101101:	sigmoid_prime = 18'b000000000000101011;
		14'b01000101101110:	sigmoid_prime = 18'b000000000000101011;
		14'b01000101101111:	sigmoid_prime = 18'b000000000000101010;
		14'b01000101110000:	sigmoid_prime = 18'b000000000000101010;
		14'b01000101110001:	sigmoid_prime = 18'b000000000000101010;
		14'b01000101110010:	sigmoid_prime = 18'b000000000000101010;
		14'b01000101110011:	sigmoid_prime = 18'b000000000000101010;
		14'b01000101110100:	sigmoid_prime = 18'b000000000000101010;
		14'b01000101110101:	sigmoid_prime = 18'b000000000000101010;
		14'b01000101110110:	sigmoid_prime = 18'b000000000000101010;
		14'b01000101110111:	sigmoid_prime = 18'b000000000000101010;
		14'b01000101111000:	sigmoid_prime = 18'b000000000000101010;
		14'b01000101111001:	sigmoid_prime = 18'b000000000000101010;
		14'b01000101111010:	sigmoid_prime = 18'b000000000000101010;
		14'b01000101111011:	sigmoid_prime = 18'b000000000000101001;
		14'b01000101111100:	sigmoid_prime = 18'b000000000000101001;
		14'b01000101111101:	sigmoid_prime = 18'b000000000000101001;
		14'b01000101111110:	sigmoid_prime = 18'b000000000000101001;
		14'b01000101111111:	sigmoid_prime = 18'b000000000000101001;
		14'b01000110000000:	sigmoid_prime = 18'b000000000000101001;
		14'b01000110000001:	sigmoid_prime = 18'b000000000000101001;
		14'b01000110000010:	sigmoid_prime = 18'b000000000000101001;
		14'b01000110000011:	sigmoid_prime = 18'b000000000000101001;
		14'b01000110000100:	sigmoid_prime = 18'b000000000000101001;
		14'b01000110000101:	sigmoid_prime = 18'b000000000000101001;
		14'b01000110000110:	sigmoid_prime = 18'b000000000000101001;
		14'b01000110000111:	sigmoid_prime = 18'b000000000000101000;
		14'b01000110001000:	sigmoid_prime = 18'b000000000000101000;
		14'b01000110001001:	sigmoid_prime = 18'b000000000000101000;
		14'b01000110001010:	sigmoid_prime = 18'b000000000000101000;
		14'b01000110001011:	sigmoid_prime = 18'b000000000000101000;
		14'b01000110001100:	sigmoid_prime = 18'b000000000000101000;
		14'b01000110001101:	sigmoid_prime = 18'b000000000000101000;
		14'b01000110001110:	sigmoid_prime = 18'b000000000000101000;
		14'b01000110001111:	sigmoid_prime = 18'b000000000000101000;
		14'b01000110010000:	sigmoid_prime = 18'b000000000000101000;
		14'b01000110010001:	sigmoid_prime = 18'b000000000000101000;
		14'b01000110010010:	sigmoid_prime = 18'b000000000000101000;
		14'b01000110010011:	sigmoid_prime = 18'b000000000000101000;
		14'b01000110010100:	sigmoid_prime = 18'b000000000000100111;
		14'b01000110010101:	sigmoid_prime = 18'b000000000000100111;
		14'b01000110010110:	sigmoid_prime = 18'b000000000000100111;
		14'b01000110010111:	sigmoid_prime = 18'b000000000000100111;
		14'b01000110011000:	sigmoid_prime = 18'b000000000000100111;
		14'b01000110011001:	sigmoid_prime = 18'b000000000000100111;
		14'b01000110011010:	sigmoid_prime = 18'b000000000000100111;
		14'b01000110011011:	sigmoid_prime = 18'b000000000000100111;
		14'b01000110011100:	sigmoid_prime = 18'b000000000000100111;
		14'b01000110011101:	sigmoid_prime = 18'b000000000000100111;
		14'b01000110011110:	sigmoid_prime = 18'b000000000000100111;
		14'b01000110011111:	sigmoid_prime = 18'b000000000000100111;
		14'b01000110100000:	sigmoid_prime = 18'b000000000000100111;
		14'b01000110100001:	sigmoid_prime = 18'b000000000000100110;
		14'b01000110100010:	sigmoid_prime = 18'b000000000000100110;
		14'b01000110100011:	sigmoid_prime = 18'b000000000000100110;
		14'b01000110100100:	sigmoid_prime = 18'b000000000000100110;
		14'b01000110100101:	sigmoid_prime = 18'b000000000000100110;
		14'b01000110100110:	sigmoid_prime = 18'b000000000000100110;
		14'b01000110100111:	sigmoid_prime = 18'b000000000000100110;
		14'b01000110101000:	sigmoid_prime = 18'b000000000000100110;
		14'b01000110101001:	sigmoid_prime = 18'b000000000000100110;
		14'b01000110101010:	sigmoid_prime = 18'b000000000000100110;
		14'b01000110101011:	sigmoid_prime = 18'b000000000000100110;
		14'b01000110101100:	sigmoid_prime = 18'b000000000000100110;
		14'b01000110101101:	sigmoid_prime = 18'b000000000000100110;
		14'b01000110101110:	sigmoid_prime = 18'b000000000000100101;
		14'b01000110101111:	sigmoid_prime = 18'b000000000000100101;
		14'b01000110110000:	sigmoid_prime = 18'b000000000000100101;
		14'b01000110110001:	sigmoid_prime = 18'b000000000000100101;
		14'b01000110110010:	sigmoid_prime = 18'b000000000000100101;
		14'b01000110110011:	sigmoid_prime = 18'b000000000000100101;
		14'b01000110110100:	sigmoid_prime = 18'b000000000000100101;
		14'b01000110110101:	sigmoid_prime = 18'b000000000000100101;
		14'b01000110110110:	sigmoid_prime = 18'b000000000000100101;
		14'b01000110110111:	sigmoid_prime = 18'b000000000000100101;
		14'b01000110111000:	sigmoid_prime = 18'b000000000000100101;
		14'b01000110111001:	sigmoid_prime = 18'b000000000000100101;
		14'b01000110111010:	sigmoid_prime = 18'b000000000000100101;
		14'b01000110111011:	sigmoid_prime = 18'b000000000000100101;
		14'b01000110111100:	sigmoid_prime = 18'b000000000000100100;
		14'b01000110111101:	sigmoid_prime = 18'b000000000000100100;
		14'b01000110111110:	sigmoid_prime = 18'b000000000000100100;
		14'b01000110111111:	sigmoid_prime = 18'b000000000000100100;
		14'b01000111000000:	sigmoid_prime = 18'b000000000000100100;
		14'b01000111000001:	sigmoid_prime = 18'b000000000000100100;
		14'b01000111000010:	sigmoid_prime = 18'b000000000000100100;
		14'b01000111000011:	sigmoid_prime = 18'b000000000000100100;
		14'b01000111000100:	sigmoid_prime = 18'b000000000000100100;
		14'b01000111000101:	sigmoid_prime = 18'b000000000000100100;
		14'b01000111000110:	sigmoid_prime = 18'b000000000000100100;
		14'b01000111000111:	sigmoid_prime = 18'b000000000000100100;
		14'b01000111001000:	sigmoid_prime = 18'b000000000000100100;
		14'b01000111001001:	sigmoid_prime = 18'b000000000000100100;
		14'b01000111001010:	sigmoid_prime = 18'b000000000000100011;
		14'b01000111001011:	sigmoid_prime = 18'b000000000000100011;
		14'b01000111001100:	sigmoid_prime = 18'b000000000000100011;
		14'b01000111001101:	sigmoid_prime = 18'b000000000000100011;
		14'b01000111001110:	sigmoid_prime = 18'b000000000000100011;
		14'b01000111001111:	sigmoid_prime = 18'b000000000000100011;
		14'b01000111010000:	sigmoid_prime = 18'b000000000000100011;
		14'b01000111010001:	sigmoid_prime = 18'b000000000000100011;
		14'b01000111010010:	sigmoid_prime = 18'b000000000000100011;
		14'b01000111010011:	sigmoid_prime = 18'b000000000000100011;
		14'b01000111010100:	sigmoid_prime = 18'b000000000000100011;
		14'b01000111010101:	sigmoid_prime = 18'b000000000000100011;
		14'b01000111010110:	sigmoid_prime = 18'b000000000000100011;
		14'b01000111010111:	sigmoid_prime = 18'b000000000000100011;
		14'b01000111011000:	sigmoid_prime = 18'b000000000000100010;
		14'b01000111011001:	sigmoid_prime = 18'b000000000000100010;
		14'b01000111011010:	sigmoid_prime = 18'b000000000000100010;
		14'b01000111011011:	sigmoid_prime = 18'b000000000000100010;
		14'b01000111011100:	sigmoid_prime = 18'b000000000000100010;
		14'b01000111011101:	sigmoid_prime = 18'b000000000000100010;
		14'b01000111011110:	sigmoid_prime = 18'b000000000000100010;
		14'b01000111011111:	sigmoid_prime = 18'b000000000000100010;
		14'b01000111100000:	sigmoid_prime = 18'b000000000000100010;
		14'b01000111100001:	sigmoid_prime = 18'b000000000000100010;
		14'b01000111100010:	sigmoid_prime = 18'b000000000000100010;
		14'b01000111100011:	sigmoid_prime = 18'b000000000000100010;
		14'b01000111100100:	sigmoid_prime = 18'b000000000000100010;
		14'b01000111100101:	sigmoid_prime = 18'b000000000000100010;
		14'b01000111100110:	sigmoid_prime = 18'b000000000000100010;
		14'b01000111100111:	sigmoid_prime = 18'b000000000000100001;
		14'b01000111101000:	sigmoid_prime = 18'b000000000000100001;
		14'b01000111101001:	sigmoid_prime = 18'b000000000000100001;
		14'b01000111101010:	sigmoid_prime = 18'b000000000000100001;
		14'b01000111101011:	sigmoid_prime = 18'b000000000000100001;
		14'b01000111101100:	sigmoid_prime = 18'b000000000000100001;
		14'b01000111101101:	sigmoid_prime = 18'b000000000000100001;
		14'b01000111101110:	sigmoid_prime = 18'b000000000000100001;
		14'b01000111101111:	sigmoid_prime = 18'b000000000000100001;
		14'b01000111110000:	sigmoid_prime = 18'b000000000000100001;
		14'b01000111110001:	sigmoid_prime = 18'b000000000000100001;
		14'b01000111110010:	sigmoid_prime = 18'b000000000000100001;
		14'b01000111110011:	sigmoid_prime = 18'b000000000000100001;
		14'b01000111110100:	sigmoid_prime = 18'b000000000000100001;
		14'b01000111110101:	sigmoid_prime = 18'b000000000000100001;
		14'b01000111110110:	sigmoid_prime = 18'b000000000000100000;
		14'b01000111110111:	sigmoid_prime = 18'b000000000000100000;
		14'b01000111111000:	sigmoid_prime = 18'b000000000000100000;
		14'b01000111111001:	sigmoid_prime = 18'b000000000000100000;
		14'b01000111111010:	sigmoid_prime = 18'b000000000000100000;
		14'b01000111111011:	sigmoid_prime = 18'b000000000000100000;
		14'b01000111111100:	sigmoid_prime = 18'b000000000000100000;
		14'b01000111111101:	sigmoid_prime = 18'b000000000000100000;
		14'b01000111111110:	sigmoid_prime = 18'b000000000000100000;
		14'b01000111111111:	sigmoid_prime = 18'b000000000000100000;
		14'b01001000000000:	sigmoid_prime = 18'b000000000000100000;
		14'b01001000000001:	sigmoid_prime = 18'b000000000000100000;
		14'b01001000000010:	sigmoid_prime = 18'b000000000000100000;
		14'b01001000000011:	sigmoid_prime = 18'b000000000000100000;
		14'b01001000000100:	sigmoid_prime = 18'b000000000000100000;
		14'b01001000000101:	sigmoid_prime = 18'b000000000000100000;
		14'b01001000000110:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000000111:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000001000:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000001001:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000001010:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000001011:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000001100:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000001101:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000001110:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000001111:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000010000:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000010001:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000010010:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000010011:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000010100:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000010101:	sigmoid_prime = 18'b000000000000011111;
		14'b01001000010110:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000010111:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000011000:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000011001:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000011010:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000011011:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000011100:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000011101:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000011110:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000011111:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000100000:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000100001:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000100010:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000100011:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000100100:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000100101:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000100110:	sigmoid_prime = 18'b000000000000011110;
		14'b01001000100111:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000101000:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000101001:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000101010:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000101011:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000101100:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000101101:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000101110:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000101111:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000110000:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000110001:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000110010:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000110011:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000110100:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000110101:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000110110:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000110111:	sigmoid_prime = 18'b000000000000011101;
		14'b01001000111000:	sigmoid_prime = 18'b000000000000011100;
		14'b01001000111001:	sigmoid_prime = 18'b000000000000011100;
		14'b01001000111010:	sigmoid_prime = 18'b000000000000011100;
		14'b01001000111011:	sigmoid_prime = 18'b000000000000011100;
		14'b01001000111100:	sigmoid_prime = 18'b000000000000011100;
		14'b01001000111101:	sigmoid_prime = 18'b000000000000011100;
		14'b01001000111110:	sigmoid_prime = 18'b000000000000011100;
		14'b01001000111111:	sigmoid_prime = 18'b000000000000011100;
		14'b01001001000000:	sigmoid_prime = 18'b000000000000011100;
		14'b01001001000001:	sigmoid_prime = 18'b000000000000011100;
		14'b01001001000010:	sigmoid_prime = 18'b000000000000011100;
		14'b01001001000011:	sigmoid_prime = 18'b000000000000011100;
		14'b01001001000100:	sigmoid_prime = 18'b000000000000011100;
		14'b01001001000101:	sigmoid_prime = 18'b000000000000011100;
		14'b01001001000110:	sigmoid_prime = 18'b000000000000011100;
		14'b01001001000111:	sigmoid_prime = 18'b000000000000011100;
		14'b01001001001000:	sigmoid_prime = 18'b000000000000011100;
		14'b01001001001001:	sigmoid_prime = 18'b000000000000011100;
		14'b01001001001010:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001001011:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001001100:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001001101:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001001110:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001001111:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001010000:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001010001:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001010010:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001010011:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001010100:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001010101:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001010110:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001010111:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001011000:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001011001:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001011010:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001011011:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001011100:	sigmoid_prime = 18'b000000000000011011;
		14'b01001001011101:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001011110:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001011111:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001100000:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001100001:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001100010:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001100011:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001100100:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001100101:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001100110:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001100111:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001101000:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001101001:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001101010:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001101011:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001101100:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001101101:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001101110:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001101111:	sigmoid_prime = 18'b000000000000011010;
		14'b01001001110000:	sigmoid_prime = 18'b000000000000011001;
		14'b01001001110001:	sigmoid_prime = 18'b000000000000011001;
		14'b01001001110010:	sigmoid_prime = 18'b000000000000011001;
		14'b01001001110011:	sigmoid_prime = 18'b000000000000011001;
		14'b01001001110100:	sigmoid_prime = 18'b000000000000011001;
		14'b01001001110101:	sigmoid_prime = 18'b000000000000011001;
		14'b01001001110110:	sigmoid_prime = 18'b000000000000011001;
		14'b01001001110111:	sigmoid_prime = 18'b000000000000011001;
		14'b01001001111000:	sigmoid_prime = 18'b000000000000011001;
		14'b01001001111001:	sigmoid_prime = 18'b000000000000011001;
		14'b01001001111010:	sigmoid_prime = 18'b000000000000011001;
		14'b01001001111011:	sigmoid_prime = 18'b000000000000011001;
		14'b01001001111100:	sigmoid_prime = 18'b000000000000011001;
		14'b01001001111101:	sigmoid_prime = 18'b000000000000011001;
		14'b01001001111110:	sigmoid_prime = 18'b000000000000011001;
		14'b01001001111111:	sigmoid_prime = 18'b000000000000011001;
		14'b01001010000000:	sigmoid_prime = 18'b000000000000011001;
		14'b01001010000001:	sigmoid_prime = 18'b000000000000011001;
		14'b01001010000010:	sigmoid_prime = 18'b000000000000011001;
		14'b01001010000011:	sigmoid_prime = 18'b000000000000011001;
		14'b01001010000100:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010000101:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010000110:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010000111:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010001000:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010001001:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010001010:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010001011:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010001100:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010001101:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010001110:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010001111:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010010000:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010010001:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010010010:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010010011:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010010100:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010010101:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010010110:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010010111:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010011000:	sigmoid_prime = 18'b000000000000011000;
		14'b01001010011001:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010011010:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010011011:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010011100:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010011101:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010011110:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010011111:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010100000:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010100001:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010100010:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010100011:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010100100:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010100101:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010100110:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010100111:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010101000:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010101001:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010101010:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010101011:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010101100:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010101101:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010101110:	sigmoid_prime = 18'b000000000000010111;
		14'b01001010101111:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010110000:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010110001:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010110010:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010110011:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010110100:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010110101:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010110110:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010110111:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010111000:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010111001:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010111010:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010111011:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010111100:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010111101:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010111110:	sigmoid_prime = 18'b000000000000010110;
		14'b01001010111111:	sigmoid_prime = 18'b000000000000010110;
		14'b01001011000000:	sigmoid_prime = 18'b000000000000010110;
		14'b01001011000001:	sigmoid_prime = 18'b000000000000010110;
		14'b01001011000010:	sigmoid_prime = 18'b000000000000010110;
		14'b01001011000011:	sigmoid_prime = 18'b000000000000010110;
		14'b01001011000100:	sigmoid_prime = 18'b000000000000010110;
		14'b01001011000101:	sigmoid_prime = 18'b000000000000010110;
		14'b01001011000110:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011000111:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011001000:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011001001:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011001010:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011001011:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011001100:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011001101:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011001110:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011001111:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011010000:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011010001:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011010010:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011010011:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011010100:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011010101:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011010110:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011010111:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011011000:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011011001:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011011010:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011011011:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011011100:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011011101:	sigmoid_prime = 18'b000000000000010101;
		14'b01001011011110:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011011111:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011100000:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011100001:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011100010:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011100011:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011100100:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011100101:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011100110:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011100111:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011101000:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011101001:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011101010:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011101011:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011101100:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011101101:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011101110:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011101111:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011110000:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011110001:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011110010:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011110011:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011110100:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011110101:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011110110:	sigmoid_prime = 18'b000000000000010100;
		14'b01001011110111:	sigmoid_prime = 18'b000000000000010011;
		14'b01001011111000:	sigmoid_prime = 18'b000000000000010011;
		14'b01001011111001:	sigmoid_prime = 18'b000000000000010011;
		14'b01001011111010:	sigmoid_prime = 18'b000000000000010011;
		14'b01001011111011:	sigmoid_prime = 18'b000000000000010011;
		14'b01001011111100:	sigmoid_prime = 18'b000000000000010011;
		14'b01001011111101:	sigmoid_prime = 18'b000000000000010011;
		14'b01001011111110:	sigmoid_prime = 18'b000000000000010011;
		14'b01001011111111:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100000000:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100000001:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100000010:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100000011:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100000100:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100000101:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100000110:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100000111:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100001000:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100001001:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100001010:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100001011:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100001100:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100001101:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100001110:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100001111:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100010000:	sigmoid_prime = 18'b000000000000010011;
		14'b01001100010001:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100010010:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100010011:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100010100:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100010101:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100010110:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100010111:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100011000:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100011001:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100011010:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100011011:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100011100:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100011101:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100011110:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100011111:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100100000:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100100001:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100100010:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100100011:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100100100:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100100101:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100100110:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100100111:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100101000:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100101001:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100101010:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100101011:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100101100:	sigmoid_prime = 18'b000000000000010010;
		14'b01001100101101:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100101110:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100101111:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100110000:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100110001:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100110010:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100110011:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100110100:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100110101:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100110110:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100110111:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100111000:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100111001:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100111010:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100111011:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100111100:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100111101:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100111110:	sigmoid_prime = 18'b000000000000010001;
		14'b01001100111111:	sigmoid_prime = 18'b000000000000010001;
		14'b01001101000000:	sigmoid_prime = 18'b000000000000010001;
		14'b01001101000001:	sigmoid_prime = 18'b000000000000010001;
		14'b01001101000010:	sigmoid_prime = 18'b000000000000010001;
		14'b01001101000011:	sigmoid_prime = 18'b000000000000010001;
		14'b01001101000100:	sigmoid_prime = 18'b000000000000010001;
		14'b01001101000101:	sigmoid_prime = 18'b000000000000010001;
		14'b01001101000110:	sigmoid_prime = 18'b000000000000010001;
		14'b01001101000111:	sigmoid_prime = 18'b000000000000010001;
		14'b01001101001000:	sigmoid_prime = 18'b000000000000010001;
		14'b01001101001001:	sigmoid_prime = 18'b000000000000010001;
		14'b01001101001010:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101001011:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101001100:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101001101:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101001110:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101001111:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101010000:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101010001:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101010010:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101010011:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101010100:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101010101:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101010110:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101010111:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101011000:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101011001:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101011010:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101011011:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101011100:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101011101:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101011110:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101011111:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101100000:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101100001:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101100010:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101100011:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101100100:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101100101:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101100110:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101100111:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101101000:	sigmoid_prime = 18'b000000000000010000;
		14'b01001101101001:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101101010:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101101011:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101101100:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101101101:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101101110:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101101111:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101110000:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101110001:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101110010:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101110011:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101110100:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101110101:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101110110:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101110111:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101111000:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101111001:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101111010:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101111011:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101111100:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101111101:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101111110:	sigmoid_prime = 18'b000000000000001111;
		14'b01001101111111:	sigmoid_prime = 18'b000000000000001111;
		14'b01001110000000:	sigmoid_prime = 18'b000000000000001111;
		14'b01001110000001:	sigmoid_prime = 18'b000000000000001111;
		14'b01001110000010:	sigmoid_prime = 18'b000000000000001111;
		14'b01001110000011:	sigmoid_prime = 18'b000000000000001111;
		14'b01001110000100:	sigmoid_prime = 18'b000000000000001111;
		14'b01001110000101:	sigmoid_prime = 18'b000000000000001111;
		14'b01001110000110:	sigmoid_prime = 18'b000000000000001111;
		14'b01001110000111:	sigmoid_prime = 18'b000000000000001111;
		14'b01001110001000:	sigmoid_prime = 18'b000000000000001111;
		14'b01001110001001:	sigmoid_prime = 18'b000000000000001111;
		14'b01001110001010:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110001011:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110001100:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110001101:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110001110:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110001111:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110010000:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110010001:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110010010:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110010011:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110010100:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110010101:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110010110:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110010111:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110011000:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110011001:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110011010:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110011011:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110011100:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110011101:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110011110:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110011111:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110100000:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110100001:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110100010:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110100011:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110100100:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110100101:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110100110:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110100111:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110101000:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110101001:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110101010:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110101011:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110101100:	sigmoid_prime = 18'b000000000000001110;
		14'b01001110101101:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110101110:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110101111:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110110000:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110110001:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110110010:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110110011:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110110100:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110110101:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110110110:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110110111:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110111000:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110111001:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110111010:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110111011:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110111100:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110111101:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110111110:	sigmoid_prime = 18'b000000000000001101;
		14'b01001110111111:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111000000:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111000001:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111000010:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111000011:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111000100:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111000101:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111000110:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111000111:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111001000:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111001001:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111001010:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111001011:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111001100:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111001101:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111001110:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111001111:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111010000:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111010001:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111010010:	sigmoid_prime = 18'b000000000000001101;
		14'b01001111010011:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111010100:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111010101:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111010110:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111010111:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111011000:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111011001:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111011010:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111011011:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111011100:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111011101:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111011110:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111011111:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111100000:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111100001:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111100010:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111100011:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111100100:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111100101:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111100110:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111100111:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111101000:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111101001:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111101010:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111101011:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111101100:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111101101:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111101110:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111101111:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111110000:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111110001:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111110010:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111110011:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111110100:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111110101:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111110110:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111110111:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111111000:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111111001:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111111010:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111111011:	sigmoid_prime = 18'b000000000000001100;
		14'b01001111111100:	sigmoid_prime = 18'b000000000000001011;
		14'b01001111111101:	sigmoid_prime = 18'b000000000000001011;
		14'b01001111111110:	sigmoid_prime = 18'b000000000000001011;
		14'b01001111111111:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000000000:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000000001:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000000010:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000000011:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000000100:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000000101:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000000110:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000000111:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000001000:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000001001:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000001010:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000001011:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000001100:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000001101:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000001110:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000001111:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000010000:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000010001:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000010010:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000010011:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000010100:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000010101:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000010110:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000010111:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000011000:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000011001:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000011010:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000011011:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000011100:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000011101:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000011110:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000011111:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000100000:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000100001:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000100010:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000100011:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000100100:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000100101:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000100110:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000100111:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000101000:	sigmoid_prime = 18'b000000000000001011;
		14'b01010000101001:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000101010:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000101011:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000101100:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000101101:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000101110:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000101111:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000110000:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000110001:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000110010:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000110011:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000110100:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000110101:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000110110:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000110111:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000111000:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000111001:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000111010:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000111011:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000111100:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000111101:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000111110:	sigmoid_prime = 18'b000000000000001010;
		14'b01010000111111:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001000000:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001000001:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001000010:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001000011:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001000100:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001000101:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001000110:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001000111:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001001000:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001001001:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001001010:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001001011:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001001100:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001001101:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001001110:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001001111:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001010000:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001010001:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001010010:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001010011:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001010100:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001010101:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001010110:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001010111:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001011000:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001011001:	sigmoid_prime = 18'b000000000000001010;
		14'b01010001011010:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001011011:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001011100:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001011101:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001011110:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001011111:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001100000:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001100001:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001100010:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001100011:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001100100:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001100101:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001100110:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001100111:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001101000:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001101001:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001101010:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001101011:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001101100:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001101101:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001101110:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001101111:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001110000:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001110001:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001110010:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001110011:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001110100:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001110101:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001110110:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001110111:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001111000:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001111001:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001111010:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001111011:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001111100:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001111101:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001111110:	sigmoid_prime = 18'b000000000000001001;
		14'b01010001111111:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010000000:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010000001:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010000010:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010000011:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010000100:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010000101:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010000110:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010000111:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010001000:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010001001:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010001010:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010001011:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010001100:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010001101:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010001110:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010001111:	sigmoid_prime = 18'b000000000000001001;
		14'b01010010010000:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010010001:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010010010:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010010011:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010010100:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010010101:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010010110:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010010111:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010011000:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010011001:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010011010:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010011011:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010011100:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010011101:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010011110:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010011111:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010100000:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010100001:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010100010:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010100011:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010100100:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010100101:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010100110:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010100111:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010101000:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010101001:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010101010:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010101011:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010101100:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010101101:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010101110:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010101111:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010110000:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010110001:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010110010:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010110011:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010110100:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010110101:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010110110:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010110111:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010111000:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010111001:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010111010:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010111011:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010111100:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010111101:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010111110:	sigmoid_prime = 18'b000000000000001000;
		14'b01010010111111:	sigmoid_prime = 18'b000000000000001000;
		14'b01010011000000:	sigmoid_prime = 18'b000000000000001000;
		14'b01010011000001:	sigmoid_prime = 18'b000000000000001000;
		14'b01010011000010:	sigmoid_prime = 18'b000000000000001000;
		14'b01010011000011:	sigmoid_prime = 18'b000000000000001000;
		14'b01010011000100:	sigmoid_prime = 18'b000000000000001000;
		14'b01010011000101:	sigmoid_prime = 18'b000000000000001000;
		14'b01010011000110:	sigmoid_prime = 18'b000000000000001000;
		14'b01010011000111:	sigmoid_prime = 18'b000000000000001000;
		14'b01010011001000:	sigmoid_prime = 18'b000000000000001000;
		14'b01010011001001:	sigmoid_prime = 18'b000000000000001000;
		14'b01010011001010:	sigmoid_prime = 18'b000000000000001000;
		14'b01010011001011:	sigmoid_prime = 18'b000000000000001000;
		14'b01010011001100:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011001101:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011001110:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011001111:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011010000:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011010001:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011010010:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011010011:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011010100:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011010101:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011010110:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011010111:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011011000:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011011001:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011011010:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011011011:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011011100:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011011101:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011011110:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011011111:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011100000:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011100001:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011100010:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011100011:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011100100:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011100101:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011100110:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011100111:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011101000:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011101001:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011101010:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011101011:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011101100:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011101101:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011101110:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011101111:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011110000:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011110001:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011110010:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011110011:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011110100:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011110101:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011110110:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011110111:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011111000:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011111001:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011111010:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011111011:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011111100:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011111101:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011111110:	sigmoid_prime = 18'b000000000000000111;
		14'b01010011111111:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100000000:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100000001:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100000010:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100000011:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100000100:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100000101:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100000110:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100000111:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100001000:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100001001:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100001010:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100001011:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100001100:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100001101:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100001110:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100001111:	sigmoid_prime = 18'b000000000000000111;
		14'b01010100010000:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100010001:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100010010:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100010011:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100010100:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100010101:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100010110:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100010111:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100011000:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100011001:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100011010:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100011011:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100011100:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100011101:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100011110:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100011111:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100100000:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100100001:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100100010:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100100011:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100100100:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100100101:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100100110:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100100111:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100101000:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100101001:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100101010:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100101011:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100101100:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100101101:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100101110:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100101111:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100110000:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100110001:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100110010:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100110011:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100110100:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100110101:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100110110:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100110111:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100111000:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100111001:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100111010:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100111011:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100111100:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100111101:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100111110:	sigmoid_prime = 18'b000000000000000110;
		14'b01010100111111:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101000000:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101000001:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101000010:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101000011:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101000100:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101000101:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101000110:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101000111:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101001000:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101001001:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101001010:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101001011:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101001100:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101001101:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101001110:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101001111:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101010000:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101010001:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101010010:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101010011:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101010100:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101010101:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101010110:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101010111:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101011000:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101011001:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101011010:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101011011:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101011100:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101011101:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101011110:	sigmoid_prime = 18'b000000000000000110;
		14'b01010101011111:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101100000:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101100001:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101100010:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101100011:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101100100:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101100101:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101100110:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101100111:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101101000:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101101001:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101101010:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101101011:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101101100:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101101101:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101101110:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101101111:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101110000:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101110001:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101110010:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101110011:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101110100:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101110101:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101110110:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101110111:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101111000:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101111001:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101111010:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101111011:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101111100:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101111101:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101111110:	sigmoid_prime = 18'b000000000000000101;
		14'b01010101111111:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110000000:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110000001:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110000010:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110000011:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110000100:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110000101:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110000110:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110000111:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110001000:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110001001:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110001010:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110001011:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110001100:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110001101:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110001110:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110001111:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110010000:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110010001:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110010010:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110010011:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110010100:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110010101:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110010110:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110010111:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110011000:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110011001:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110011010:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110011011:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110011100:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110011101:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110011110:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110011111:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110100000:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110100001:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110100010:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110100011:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110100100:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110100101:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110100110:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110100111:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110101000:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110101001:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110101010:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110101011:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110101100:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110101101:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110101110:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110101111:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110110000:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110110001:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110110010:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110110011:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110110100:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110110101:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110110110:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110110111:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110111000:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110111001:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110111010:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110111011:	sigmoid_prime = 18'b000000000000000101;
		14'b01010110111100:	sigmoid_prime = 18'b000000000000000100;
		14'b01010110111101:	sigmoid_prime = 18'b000000000000000100;
		14'b01010110111110:	sigmoid_prime = 18'b000000000000000100;
		14'b01010110111111:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111000000:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111000001:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111000010:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111000011:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111000100:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111000101:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111000110:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111000111:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111001000:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111001001:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111001010:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111001011:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111001100:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111001101:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111001110:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111001111:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111010000:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111010001:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111010010:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111010011:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111010100:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111010101:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111010110:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111010111:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111011000:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111011001:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111011010:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111011011:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111011100:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111011101:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111011110:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111011111:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111100000:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111100001:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111100010:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111100011:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111100100:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111100101:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111100110:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111100111:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111101000:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111101001:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111101010:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111101011:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111101100:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111101101:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111101110:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111101111:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111110000:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111110001:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111110010:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111110011:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111110100:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111110101:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111110110:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111110111:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111111000:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111111001:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111111010:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111111011:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111111100:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111111101:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111111110:	sigmoid_prime = 18'b000000000000000100;
		14'b01010111111111:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000000000:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000000001:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000000010:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000000011:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000000100:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000000101:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000000110:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000000111:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000001000:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000001001:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000001010:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000001011:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000001100:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000001101:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000001110:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000001111:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000010000:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000010001:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000010010:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000010011:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000010100:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000010101:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000010110:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000010111:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000011000:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000011001:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000011010:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000011011:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000011100:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000011101:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000011110:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000011111:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000100000:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000100001:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000100010:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000100011:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000100100:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000100101:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000100110:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000100111:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000101000:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000101001:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000101010:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000101011:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000101100:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000101101:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000101110:	sigmoid_prime = 18'b000000000000000100;
		14'b01011000101111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000110000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000110001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000110010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000110011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000110100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000110101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000110110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000110111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000111000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000111001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000111010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000111011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000111100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000111101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000111110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011000111111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001000000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001000001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001000010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001000011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001000100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001000101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001000110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001000111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001001000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001001001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001001010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001001011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001001100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001001101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001001110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001001111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001010000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001010001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001010010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001010011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001010100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001010101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001010110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001010111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001011000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001011001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001011010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001011011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001011100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001011101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001011110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001011111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001100000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001100001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001100010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001100011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001100100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001100101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001100110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001100111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001101000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001101001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001101010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001101011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001101100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001101101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001101110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001101111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001110000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001110001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001110010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001110011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001110100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001110101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001110110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001110111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001111000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001111001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001111010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001111011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001111100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001111101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001111110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011001111111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010000000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010000001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010000010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010000011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010000100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010000101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010000110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010000111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010001000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010001001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010001010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010001011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010001100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010001101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010001110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010001111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010010000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010010001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010010010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010010011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010010100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010010101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010010110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010010111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010011000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010011001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010011010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010011011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010011100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010011101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010011110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010011111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010100000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010100001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010100010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010100011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010100100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010100101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010100110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010100111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010101000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010101001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010101010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010101011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010101100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010101101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010101110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010101111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010110000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010110001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010110010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010110011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010110100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010110101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010110110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010110111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010111000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010111001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010111010:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010111011:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010111100:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010111101:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010111110:	sigmoid_prime = 18'b000000000000000011;
		14'b01011010111111:	sigmoid_prime = 18'b000000000000000011;
		14'b01011011000000:	sigmoid_prime = 18'b000000000000000011;
		14'b01011011000001:	sigmoid_prime = 18'b000000000000000011;
		14'b01011011000010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011000011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011000100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011000101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011000110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011000111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011001000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011001001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011001010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011001011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011001100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011001101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011001110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011001111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011010000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011010001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011010010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011010011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011010100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011010101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011010110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011010111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011011000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011011001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011011010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011011011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011011100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011011101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011011110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011011111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011100000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011100001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011100010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011100011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011100100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011100101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011100110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011100111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011101000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011101001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011101010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011101011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011101100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011101101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011101110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011101111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011110000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011110001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011110010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011110011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011110100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011110101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011110110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011110111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011111000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011111001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011111010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011111011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011111100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011111101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011111110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011011111111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100000000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100000001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100000010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100000011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100000100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100000101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100000110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100000111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100001000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100001001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100001010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100001011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100001100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100001101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100001110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100001111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100010000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100010001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100010010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100010011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100010100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100010101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100010110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100010111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100011000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100011001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100011010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100011011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100011100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100011101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100011110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100011111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100100000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100100001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100100010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100100011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100100100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100100101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100100110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100100111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100101000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100101001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100101010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100101011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100101100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100101101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100101110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100101111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100110000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100110001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100110010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100110011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100110100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100110101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100110110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100110111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100111000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100111001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100111010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100111011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100111100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100111101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100111110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011100111111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101000000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101000001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101000010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101000011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101000100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101000101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101000110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101000111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101001000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101001001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101001010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101001011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101001100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101001101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101001110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101001111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101010000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101010001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101010010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101010011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101010100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101010101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101010110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101010111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101011000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101011001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101011010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101011011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101011100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101011101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101011110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101011111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101100000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101100001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101100010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101100011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101100100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101100101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101100110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101100111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101101000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101101001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101101010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101101011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101101100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101101101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101101110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101101111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101110000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101110001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101110010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101110011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101110100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101110101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101110110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101110111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101111000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101111001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101111010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101111011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101111100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101111101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101111110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011101111111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110000000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110000001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110000010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110000011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110000100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110000101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110000110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110000111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110001000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110001001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110001010:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110001011:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110001100:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110001101:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110001110:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110001111:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110010000:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110010001:	sigmoid_prime = 18'b000000000000000010;
		14'b01011110010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01011110111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01011111111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100000111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100001111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100010111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100011111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100100111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100101111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100110111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01100111111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101000111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101001111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101010111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101011111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101100111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101101111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101110111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01101111111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110000111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110001111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110010111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110011111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110100111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110101111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110110111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01110111111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111000111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111001111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111010111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111011111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111100111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111101111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111110111111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111000000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111000001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111000010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111000011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111000100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111000101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111000110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111000111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111001000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111001001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111001010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111001011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111001100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111001101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111001110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111001111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111010000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111010001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111010010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111010011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111010100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111010101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111010110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111010111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111011000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111011001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111011010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111011011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111011100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111011101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111011110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111011111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111100000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111100001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111100010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111100011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111100100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111100101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111100110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111100111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111101000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111101001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111101010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111101011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111101100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111101101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111101110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111101111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111110000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111110001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111110010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111110011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111110100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111110101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111110110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111110111:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111111000:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111111001:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111111010:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111111011:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111111100:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111111101:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111111110:	sigmoid_prime = 18'b000000000000000001;
		14'b01111111111111:	sigmoid_prime = 18'b000000000000000001;


	endcase
endmodule
