// If any parameter is changed, tables will have to be regenerated using dnn-rtl/scripts/actlut_generator.py
// TO BE REPLACED: parameter values, and the table portion inside the case statements
// NOTHING ELSE NEEDS TO BE REPLACED APART FROM ABOVE

`timescale 1ns/100ps

module sigmoid_t #(
	parameter width = 10,
	parameter int_bits = 2,
	parameter frac_bits = width-int_bits-1,
	parameter maxdomain = (2**int_bits>8) ? 8 : 2**int_bits, //8 is arbitrarily chosen
	//input has to be within [-maxdomain,maxdomain). If outside this range, sigmoid is either 0 or 1
	parameter lut_size = (2**width>4096) ? 4096 : 2**width //no. of cells in LUT
)(
	input clk,
	input signed [width-1:0] z,
	output reg [width-1:0] sigmoid_out
);
	reg [frac_bits-1:0] sigmoid;

	/*always @(posedge clk)
		if(z[width-1]==1|| z==0 )
			sigmoid_out = (z[width-1:width-int_bits+2] == 0 || (&z[width-1:width-int_bits+2] ))?
			{{(int_bits+1){1'b0}}, sigmoid}: 
			(z[width-1])?  1: {1'b1, {(frac_bits){1'b0}}}-1;
		else
			sigmoid_out = z;*/

	always @(posedge clk) begin
		sigmoid_out = (z[width-1:width-int_bits+$clog2(maxdomain)-1] == 0 || &z[width-1:width-int_bits+$clog2(maxdomain)-1]) ? // Only calculate sigmoid for the domain z = [-maxdomain,+maxdomain). So check all MSB till there. If all 0, z<8. If all 1, z>=-8
		{{(int_bits+1){1'b0}}, sigmoid} : //If z is within [-maxdomain,+maxdomain), insert all 0s for sign and integer part (since sigmoid is always between 0 and 1) and then frac_bits sigmoid part
		(z[width-1]) ? //If z is outside the range, sigmoid will be 0 or 1 depending on sign bit
		1 : //If sign bit is 1, z is negative. Then sigmoid is all zeros followed by 1 at LSB, i.e. 2^(-frac_bits), which is the lowest number possible (~=0)
		{{(int_bits+1){1'b0}},{(frac_bits){1'b1}}}; //If sign bit is 0, z is positive. Then sigmoid is all 1s in the frational part, i.e. 1-2^(-frac_bits), which is the highest number possible (~=1)
	end

	always @(z[frac_bits+$clog2(maxdomain):frac_bits-$clog2(lut_size)+$clog2(maxdomain)+1]) //this ensures that we read exactly log(lut_size) bits as address of LUT
	case (z[frac_bits+$clog2(maxdomain):frac_bits-$clog2(lut_size)+$clog2(maxdomain)+1])

		10'b1000000000:	sigmoid = 7'b0000010;
		10'b1000000001:	sigmoid = 7'b0000010;
		10'b1000000010:	sigmoid = 7'b0000010;
		10'b1000000011:	sigmoid = 7'b0000010;
		10'b1000000100:	sigmoid = 7'b0000010;
		10'b1000000101:	sigmoid = 7'b0000010;
		10'b1000000110:	sigmoid = 7'b0000010;
		10'b1000000111:	sigmoid = 7'b0000010;
		10'b1000001000:	sigmoid = 7'b0000010;
		10'b1000001001:	sigmoid = 7'b0000010;
		10'b1000001010:	sigmoid = 7'b0000010;
		10'b1000001011:	sigmoid = 7'b0000011;
		10'b1000001100:	sigmoid = 7'b0000011;
		10'b1000001101:	sigmoid = 7'b0000011;
		10'b1000001110:	sigmoid = 7'b0000011;
		10'b1000001111:	sigmoid = 7'b0000011;
		10'b1000010000:	sigmoid = 7'b0000011;
		10'b1000010001:	sigmoid = 7'b0000011;
		10'b1000010010:	sigmoid = 7'b0000011;
		10'b1000010011:	sigmoid = 7'b0000011;
		10'b1000010100:	sigmoid = 7'b0000011;
		10'b1000010101:	sigmoid = 7'b0000011;
		10'b1000010110:	sigmoid = 7'b0000011;
		10'b1000010111:	sigmoid = 7'b0000011;
		10'b1000011000:	sigmoid = 7'b0000011;
		10'b1000011001:	sigmoid = 7'b0000011;
		10'b1000011010:	sigmoid = 7'b0000011;
		10'b1000011011:	sigmoid = 7'b0000011;
		10'b1000011100:	sigmoid = 7'b0000011;
		10'b1000011101:	sigmoid = 7'b0000011;
		10'b1000011110:	sigmoid = 7'b0000011;
		10'b1000011111:	sigmoid = 7'b0000011;
		10'b1000100000:	sigmoid = 7'b0000011;
		10'b1000100001:	sigmoid = 7'b0000011;
		10'b1000100010:	sigmoid = 7'b0000011;
		10'b1000100011:	sigmoid = 7'b0000011;
		10'b1000100100:	sigmoid = 7'b0000011;
		10'b1000100101:	sigmoid = 7'b0000011;
		10'b1000100110:	sigmoid = 7'b0000011;
		10'b1000100111:	sigmoid = 7'b0000011;
		10'b1000101000:	sigmoid = 7'b0000011;
		10'b1000101001:	sigmoid = 7'b0000011;
		10'b1000101010:	sigmoid = 7'b0000011;
		10'b1000101011:	sigmoid = 7'b0000011;
		10'b1000101100:	sigmoid = 7'b0000011;
		10'b1000101101:	sigmoid = 7'b0000011;
		10'b1000101110:	sigmoid = 7'b0000011;
		10'b1000101111:	sigmoid = 7'b0000011;
		10'b1000110000:	sigmoid = 7'b0000011;
		10'b1000110001:	sigmoid = 7'b0000011;
		10'b1000110010:	sigmoid = 7'b0000011;
		10'b1000110011:	sigmoid = 7'b0000011;
		10'b1000110100:	sigmoid = 7'b0000011;
		10'b1000110101:	sigmoid = 7'b0000011;
		10'b1000110110:	sigmoid = 7'b0000011;
		10'b1000110111:	sigmoid = 7'b0000100;
		10'b1000111000:	sigmoid = 7'b0000100;
		10'b1000111001:	sigmoid = 7'b0000100;
		10'b1000111010:	sigmoid = 7'b0000100;
		10'b1000111011:	sigmoid = 7'b0000100;
		10'b1000111100:	sigmoid = 7'b0000100;
		10'b1000111101:	sigmoid = 7'b0000100;
		10'b1000111110:	sigmoid = 7'b0000100;
		10'b1000111111:	sigmoid = 7'b0000100;
		10'b1001000000:	sigmoid = 7'b0000100;
		10'b1001000001:	sigmoid = 7'b0000100;
		10'b1001000010:	sigmoid = 7'b0000100;
		10'b1001000011:	sigmoid = 7'b0000100;
		10'b1001000100:	sigmoid = 7'b0000100;
		10'b1001000101:	sigmoid = 7'b0000100;
		10'b1001000110:	sigmoid = 7'b0000100;
		10'b1001000111:	sigmoid = 7'b0000100;
		10'b1001001000:	sigmoid = 7'b0000100;
		10'b1001001001:	sigmoid = 7'b0000100;
		10'b1001001010:	sigmoid = 7'b0000100;
		10'b1001001011:	sigmoid = 7'b0000100;
		10'b1001001100:	sigmoid = 7'b0000100;
		10'b1001001101:	sigmoid = 7'b0000100;
		10'b1001001110:	sigmoid = 7'b0000100;
		10'b1001001111:	sigmoid = 7'b0000100;
		10'b1001010000:	sigmoid = 7'b0000100;
		10'b1001010001:	sigmoid = 7'b0000100;
		10'b1001010010:	sigmoid = 7'b0000100;
		10'b1001010011:	sigmoid = 7'b0000100;
		10'b1001010100:	sigmoid = 7'b0000100;
		10'b1001010101:	sigmoid = 7'b0000100;
		10'b1001010110:	sigmoid = 7'b0000100;
		10'b1001010111:	sigmoid = 7'b0000100;
		10'b1001011000:	sigmoid = 7'b0000100;
		10'b1001011001:	sigmoid = 7'b0000101;
		10'b1001011010:	sigmoid = 7'b0000101;
		10'b1001011011:	sigmoid = 7'b0000101;
		10'b1001011100:	sigmoid = 7'b0000101;
		10'b1001011101:	sigmoid = 7'b0000101;
		10'b1001011110:	sigmoid = 7'b0000101;
		10'b1001011111:	sigmoid = 7'b0000101;
		10'b1001100000:	sigmoid = 7'b0000101;
		10'b1001100001:	sigmoid = 7'b0000101;
		10'b1001100010:	sigmoid = 7'b0000101;
		10'b1001100011:	sigmoid = 7'b0000101;
		10'b1001100100:	sigmoid = 7'b0000101;
		10'b1001100101:	sigmoid = 7'b0000101;
		10'b1001100110:	sigmoid = 7'b0000101;
		10'b1001100111:	sigmoid = 7'b0000101;
		10'b1001101000:	sigmoid = 7'b0000101;
		10'b1001101001:	sigmoid = 7'b0000101;
		10'b1001101010:	sigmoid = 7'b0000101;
		10'b1001101011:	sigmoid = 7'b0000101;
		10'b1001101100:	sigmoid = 7'b0000101;
		10'b1001101101:	sigmoid = 7'b0000101;
		10'b1001101110:	sigmoid = 7'b0000101;
		10'b1001101111:	sigmoid = 7'b0000101;
		10'b1001110000:	sigmoid = 7'b0000101;
		10'b1001110001:	sigmoid = 7'b0000101;
		10'b1001110010:	sigmoid = 7'b0000101;
		10'b1001110011:	sigmoid = 7'b0000110;
		10'b1001110100:	sigmoid = 7'b0000110;
		10'b1001110101:	sigmoid = 7'b0000110;
		10'b1001110110:	sigmoid = 7'b0000110;
		10'b1001110111:	sigmoid = 7'b0000110;
		10'b1001111000:	sigmoid = 7'b0000110;
		10'b1001111001:	sigmoid = 7'b0000110;
		10'b1001111010:	sigmoid = 7'b0000110;
		10'b1001111011:	sigmoid = 7'b0000110;
		10'b1001111100:	sigmoid = 7'b0000110;
		10'b1001111101:	sigmoid = 7'b0000110;
		10'b1001111110:	sigmoid = 7'b0000110;
		10'b1001111111:	sigmoid = 7'b0000110;
		10'b1010000000:	sigmoid = 7'b0000110;
		10'b1010000001:	sigmoid = 7'b0000110;
		10'b1010000010:	sigmoid = 7'b0000110;
		10'b1010000011:	sigmoid = 7'b0000110;
		10'b1010000100:	sigmoid = 7'b0000110;
		10'b1010000101:	sigmoid = 7'b0000110;
		10'b1010000110:	sigmoid = 7'b0000110;
		10'b1010000111:	sigmoid = 7'b0000110;
		10'b1010001000:	sigmoid = 7'b0000110;
		10'b1010001001:	sigmoid = 7'b0000110;
		10'b1010001010:	sigmoid = 7'b0000111;
		10'b1010001011:	sigmoid = 7'b0000111;
		10'b1010001100:	sigmoid = 7'b0000111;
		10'b1010001101:	sigmoid = 7'b0000111;
		10'b1010001110:	sigmoid = 7'b0000111;
		10'b1010001111:	sigmoid = 7'b0000111;
		10'b1010010000:	sigmoid = 7'b0000111;
		10'b1010010001:	sigmoid = 7'b0000111;
		10'b1010010010:	sigmoid = 7'b0000111;
		10'b1010010011:	sigmoid = 7'b0000111;
		10'b1010010100:	sigmoid = 7'b0000111;
		10'b1010010101:	sigmoid = 7'b0000111;
		10'b1010010110:	sigmoid = 7'b0000111;
		10'b1010010111:	sigmoid = 7'b0000111;
		10'b1010011000:	sigmoid = 7'b0000111;
		10'b1010011001:	sigmoid = 7'b0000111;
		10'b1010011010:	sigmoid = 7'b0000111;
		10'b1010011011:	sigmoid = 7'b0000111;
		10'b1010011100:	sigmoid = 7'b0000111;
		10'b1010011101:	sigmoid = 7'b0001000;
		10'b1010011110:	sigmoid = 7'b0001000;
		10'b1010011111:	sigmoid = 7'b0001000;
		10'b1010100000:	sigmoid = 7'b0001000;
		10'b1010100001:	sigmoid = 7'b0001000;
		10'b1010100010:	sigmoid = 7'b0001000;
		10'b1010100011:	sigmoid = 7'b0001000;
		10'b1010100100:	sigmoid = 7'b0001000;
		10'b1010100101:	sigmoid = 7'b0001000;
		10'b1010100110:	sigmoid = 7'b0001000;
		10'b1010100111:	sigmoid = 7'b0001000;
		10'b1010101000:	sigmoid = 7'b0001000;
		10'b1010101001:	sigmoid = 7'b0001000;
		10'b1010101010:	sigmoid = 7'b0001000;
		10'b1010101011:	sigmoid = 7'b0001000;
		10'b1010101100:	sigmoid = 7'b0001000;
		10'b1010101101:	sigmoid = 7'b0001000;
		10'b1010101110:	sigmoid = 7'b0001001;
		10'b1010101111:	sigmoid = 7'b0001001;
		10'b1010110000:	sigmoid = 7'b0001001;
		10'b1010110001:	sigmoid = 7'b0001001;
		10'b1010110010:	sigmoid = 7'b0001001;
		10'b1010110011:	sigmoid = 7'b0001001;
		10'b1010110100:	sigmoid = 7'b0001001;
		10'b1010110101:	sigmoid = 7'b0001001;
		10'b1010110110:	sigmoid = 7'b0001001;
		10'b1010110111:	sigmoid = 7'b0001001;
		10'b1010111000:	sigmoid = 7'b0001001;
		10'b1010111001:	sigmoid = 7'b0001001;
		10'b1010111010:	sigmoid = 7'b0001001;
		10'b1010111011:	sigmoid = 7'b0001001;
		10'b1010111100:	sigmoid = 7'b0001001;
		10'b1010111101:	sigmoid = 7'b0001010;
		10'b1010111110:	sigmoid = 7'b0001010;
		10'b1010111111:	sigmoid = 7'b0001010;
		10'b1011000000:	sigmoid = 7'b0001010;
		10'b1011000001:	sigmoid = 7'b0001010;
		10'b1011000010:	sigmoid = 7'b0001010;
		10'b1011000011:	sigmoid = 7'b0001010;
		10'b1011000100:	sigmoid = 7'b0001010;
		10'b1011000101:	sigmoid = 7'b0001010;
		10'b1011000110:	sigmoid = 7'b0001010;
		10'b1011000111:	sigmoid = 7'b0001010;
		10'b1011001000:	sigmoid = 7'b0001010;
		10'b1011001001:	sigmoid = 7'b0001010;
		10'b1011001010:	sigmoid = 7'b0001010;
		10'b1011001011:	sigmoid = 7'b0001011;
		10'b1011001100:	sigmoid = 7'b0001011;
		10'b1011001101:	sigmoid = 7'b0001011;
		10'b1011001110:	sigmoid = 7'b0001011;
		10'b1011001111:	sigmoid = 7'b0001011;
		10'b1011010000:	sigmoid = 7'b0001011;
		10'b1011010001:	sigmoid = 7'b0001011;
		10'b1011010010:	sigmoid = 7'b0001011;
		10'b1011010011:	sigmoid = 7'b0001011;
		10'b1011010100:	sigmoid = 7'b0001011;
		10'b1011010101:	sigmoid = 7'b0001011;
		10'b1011010110:	sigmoid = 7'b0001011;
		10'b1011010111:	sigmoid = 7'b0001011;
		10'b1011011000:	sigmoid = 7'b0001100;
		10'b1011011001:	sigmoid = 7'b0001100;
		10'b1011011010:	sigmoid = 7'b0001100;
		10'b1011011011:	sigmoid = 7'b0001100;
		10'b1011011100:	sigmoid = 7'b0001100;
		10'b1011011101:	sigmoid = 7'b0001100;
		10'b1011011110:	sigmoid = 7'b0001100;
		10'b1011011111:	sigmoid = 7'b0001100;
		10'b1011100000:	sigmoid = 7'b0001100;
		10'b1011100001:	sigmoid = 7'b0001100;
		10'b1011100010:	sigmoid = 7'b0001100;
		10'b1011100011:	sigmoid = 7'b0001100;
		10'b1011100100:	sigmoid = 7'b0001101;
		10'b1011100101:	sigmoid = 7'b0001101;
		10'b1011100110:	sigmoid = 7'b0001101;
		10'b1011100111:	sigmoid = 7'b0001101;
		10'b1011101000:	sigmoid = 7'b0001101;
		10'b1011101001:	sigmoid = 7'b0001101;
		10'b1011101010:	sigmoid = 7'b0001101;
		10'b1011101011:	sigmoid = 7'b0001101;
		10'b1011101100:	sigmoid = 7'b0001101;
		10'b1011101101:	sigmoid = 7'b0001101;
		10'b1011101110:	sigmoid = 7'b0001101;
		10'b1011101111:	sigmoid = 7'b0001110;
		10'b1011110000:	sigmoid = 7'b0001110;
		10'b1011110001:	sigmoid = 7'b0001110;
		10'b1011110010:	sigmoid = 7'b0001110;
		10'b1011110011:	sigmoid = 7'b0001110;
		10'b1011110100:	sigmoid = 7'b0001110;
		10'b1011110101:	sigmoid = 7'b0001110;
		10'b1011110110:	sigmoid = 7'b0001110;
		10'b1011110111:	sigmoid = 7'b0001110;
		10'b1011111000:	sigmoid = 7'b0001110;
		10'b1011111001:	sigmoid = 7'b0001111;
		10'b1011111010:	sigmoid = 7'b0001111;
		10'b1011111011:	sigmoid = 7'b0001111;
		10'b1011111100:	sigmoid = 7'b0001111;
		10'b1011111101:	sigmoid = 7'b0001111;
		10'b1011111110:	sigmoid = 7'b0001111;
		10'b1011111111:	sigmoid = 7'b0001111;
		10'b1100000000:	sigmoid = 7'b0001111;
		10'b1100000001:	sigmoid = 7'b0001111;
		10'b1100000010:	sigmoid = 7'b0001111;
		10'b1100000011:	sigmoid = 7'b0010000;
		10'b1100000100:	sigmoid = 7'b0010000;
		10'b1100000101:	sigmoid = 7'b0010000;
		10'b1100000110:	sigmoid = 7'b0010000;
		10'b1100000111:	sigmoid = 7'b0010000;
		10'b1100001000:	sigmoid = 7'b0010000;
		10'b1100001001:	sigmoid = 7'b0010000;
		10'b1100001010:	sigmoid = 7'b0010000;
		10'b1100001011:	sigmoid = 7'b0010000;
		10'b1100001100:	sigmoid = 7'b0010001;
		10'b1100001101:	sigmoid = 7'b0010001;
		10'b1100001110:	sigmoid = 7'b0010001;
		10'b1100001111:	sigmoid = 7'b0010001;
		10'b1100010000:	sigmoid = 7'b0010001;
		10'b1100010001:	sigmoid = 7'b0010001;
		10'b1100010010:	sigmoid = 7'b0010001;
		10'b1100010011:	sigmoid = 7'b0010001;
		10'b1100010100:	sigmoid = 7'b0010001;
		10'b1100010101:	sigmoid = 7'b0010010;
		10'b1100010110:	sigmoid = 7'b0010010;
		10'b1100010111:	sigmoid = 7'b0010010;
		10'b1100011000:	sigmoid = 7'b0010010;
		10'b1100011001:	sigmoid = 7'b0010010;
		10'b1100011010:	sigmoid = 7'b0010010;
		10'b1100011011:	sigmoid = 7'b0010010;
		10'b1100011100:	sigmoid = 7'b0010010;
		10'b1100011101:	sigmoid = 7'b0010011;
		10'b1100011110:	sigmoid = 7'b0010011;
		10'b1100011111:	sigmoid = 7'b0010011;
		10'b1100100000:	sigmoid = 7'b0010011;
		10'b1100100001:	sigmoid = 7'b0010011;
		10'b1100100010:	sigmoid = 7'b0010011;
		10'b1100100011:	sigmoid = 7'b0010011;
		10'b1100100100:	sigmoid = 7'b0010011;
		10'b1100100101:	sigmoid = 7'b0010100;
		10'b1100100110:	sigmoid = 7'b0010100;
		10'b1100100111:	sigmoid = 7'b0010100;
		10'b1100101000:	sigmoid = 7'b0010100;
		10'b1100101001:	sigmoid = 7'b0010100;
		10'b1100101010:	sigmoid = 7'b0010100;
		10'b1100101011:	sigmoid = 7'b0010100;
		10'b1100101100:	sigmoid = 7'b0010101;
		10'b1100101101:	sigmoid = 7'b0010101;
		10'b1100101110:	sigmoid = 7'b0010101;
		10'b1100101111:	sigmoid = 7'b0010101;
		10'b1100110000:	sigmoid = 7'b0010101;
		10'b1100110001:	sigmoid = 7'b0010101;
		10'b1100110010:	sigmoid = 7'b0010101;
		10'b1100110011:	sigmoid = 7'b0010101;
		10'b1100110100:	sigmoid = 7'b0010110;
		10'b1100110101:	sigmoid = 7'b0010110;
		10'b1100110110:	sigmoid = 7'b0010110;
		10'b1100110111:	sigmoid = 7'b0010110;
		10'b1100111000:	sigmoid = 7'b0010110;
		10'b1100111001:	sigmoid = 7'b0010110;
		10'b1100111010:	sigmoid = 7'b0010110;
		10'b1100111011:	sigmoid = 7'b0010111;
		10'b1100111100:	sigmoid = 7'b0010111;
		10'b1100111101:	sigmoid = 7'b0010111;
		10'b1100111110:	sigmoid = 7'b0010111;
		10'b1100111111:	sigmoid = 7'b0010111;
		10'b1101000000:	sigmoid = 7'b0010111;
		10'b1101000001:	sigmoid = 7'b0010111;
		10'b1101000010:	sigmoid = 7'b0011000;
		10'b1101000011:	sigmoid = 7'b0011000;
		10'b1101000100:	sigmoid = 7'b0011000;
		10'b1101000101:	sigmoid = 7'b0011000;
		10'b1101000110:	sigmoid = 7'b0011000;
		10'b1101000111:	sigmoid = 7'b0011000;
		10'b1101001000:	sigmoid = 7'b0011001;
		10'b1101001001:	sigmoid = 7'b0011001;
		10'b1101001010:	sigmoid = 7'b0011001;
		10'b1101001011:	sigmoid = 7'b0011001;
		10'b1101001100:	sigmoid = 7'b0011001;
		10'b1101001101:	sigmoid = 7'b0011001;
		10'b1101001110:	sigmoid = 7'b0011010;
		10'b1101001111:	sigmoid = 7'b0011010;
		10'b1101010000:	sigmoid = 7'b0011010;
		10'b1101010001:	sigmoid = 7'b0011010;
		10'b1101010010:	sigmoid = 7'b0011010;
		10'b1101010011:	sigmoid = 7'b0011010;
		10'b1101010100:	sigmoid = 7'b0011010;
		10'b1101010101:	sigmoid = 7'b0011011;
		10'b1101010110:	sigmoid = 7'b0011011;
		10'b1101010111:	sigmoid = 7'b0011011;
		10'b1101011000:	sigmoid = 7'b0011011;
		10'b1101011001:	sigmoid = 7'b0011011;
		10'b1101011010:	sigmoid = 7'b0011011;
		10'b1101011011:	sigmoid = 7'b0011100;
		10'b1101011100:	sigmoid = 7'b0011100;
		10'b1101011101:	sigmoid = 7'b0011100;
		10'b1101011110:	sigmoid = 7'b0011100;
		10'b1101011111:	sigmoid = 7'b0011100;
		10'b1101100000:	sigmoid = 7'b0011101;
		10'b1101100001:	sigmoid = 7'b0011101;
		10'b1101100010:	sigmoid = 7'b0011101;
		10'b1101100011:	sigmoid = 7'b0011101;
		10'b1101100100:	sigmoid = 7'b0011101;
		10'b1101100101:	sigmoid = 7'b0011101;
		10'b1101100110:	sigmoid = 7'b0011110;
		10'b1101100111:	sigmoid = 7'b0011110;
		10'b1101101000:	sigmoid = 7'b0011110;
		10'b1101101001:	sigmoid = 7'b0011110;
		10'b1101101010:	sigmoid = 7'b0011110;
		10'b1101101011:	sigmoid = 7'b0011110;
		10'b1101101100:	sigmoid = 7'b0011111;
		10'b1101101101:	sigmoid = 7'b0011111;
		10'b1101101110:	sigmoid = 7'b0011111;
		10'b1101101111:	sigmoid = 7'b0011111;
		10'b1101110000:	sigmoid = 7'b0011111;
		10'b1101110001:	sigmoid = 7'b0100000;
		10'b1101110010:	sigmoid = 7'b0100000;
		10'b1101110011:	sigmoid = 7'b0100000;
		10'b1101110100:	sigmoid = 7'b0100000;
		10'b1101110101:	sigmoid = 7'b0100000;
		10'b1101110110:	sigmoid = 7'b0100000;
		10'b1101110111:	sigmoid = 7'b0100001;
		10'b1101111000:	sigmoid = 7'b0100001;
		10'b1101111001:	sigmoid = 7'b0100001;
		10'b1101111010:	sigmoid = 7'b0100001;
		10'b1101111011:	sigmoid = 7'b0100001;
		10'b1101111100:	sigmoid = 7'b0100010;
		10'b1101111101:	sigmoid = 7'b0100010;
		10'b1101111110:	sigmoid = 7'b0100010;
		10'b1101111111:	sigmoid = 7'b0100010;
		10'b1110000000:	sigmoid = 7'b0100010;
		10'b1110000001:	sigmoid = 7'b0100011;
		10'b1110000010:	sigmoid = 7'b0100011;
		10'b1110000011:	sigmoid = 7'b0100011;
		10'b1110000100:	sigmoid = 7'b0100011;
		10'b1110000101:	sigmoid = 7'b0100011;
		10'b1110000110:	sigmoid = 7'b0100100;
		10'b1110000111:	sigmoid = 7'b0100100;
		10'b1110001000:	sigmoid = 7'b0100100;
		10'b1110001001:	sigmoid = 7'b0100100;
		10'b1110001010:	sigmoid = 7'b0100100;
		10'b1110001011:	sigmoid = 7'b0100101;
		10'b1110001100:	sigmoid = 7'b0100101;
		10'b1110001101:	sigmoid = 7'b0100101;
		10'b1110001110:	sigmoid = 7'b0100101;
		10'b1110001111:	sigmoid = 7'b0100101;
		10'b1110010000:	sigmoid = 7'b0100110;
		10'b1110010001:	sigmoid = 7'b0100110;
		10'b1110010010:	sigmoid = 7'b0100110;
		10'b1110010011:	sigmoid = 7'b0100110;
		10'b1110010100:	sigmoid = 7'b0100110;
		10'b1110010101:	sigmoid = 7'b0100111;
		10'b1110010110:	sigmoid = 7'b0100111;
		10'b1110010111:	sigmoid = 7'b0100111;
		10'b1110011000:	sigmoid = 7'b0100111;
		10'b1110011001:	sigmoid = 7'b0101000;
		10'b1110011010:	sigmoid = 7'b0101000;
		10'b1110011011:	sigmoid = 7'b0101000;
		10'b1110011100:	sigmoid = 7'b0101000;
		10'b1110011101:	sigmoid = 7'b0101000;
		10'b1110011110:	sigmoid = 7'b0101001;
		10'b1110011111:	sigmoid = 7'b0101001;
		10'b1110100000:	sigmoid = 7'b0101001;
		10'b1110100001:	sigmoid = 7'b0101001;
		10'b1110100010:	sigmoid = 7'b0101010;
		10'b1110100011:	sigmoid = 7'b0101010;
		10'b1110100100:	sigmoid = 7'b0101010;
		10'b1110100101:	sigmoid = 7'b0101010;
		10'b1110100110:	sigmoid = 7'b0101010;
		10'b1110100111:	sigmoid = 7'b0101011;
		10'b1110101000:	sigmoid = 7'b0101011;
		10'b1110101001:	sigmoid = 7'b0101011;
		10'b1110101010:	sigmoid = 7'b0101011;
		10'b1110101011:	sigmoid = 7'b0101011;
		10'b1110101100:	sigmoid = 7'b0101100;
		10'b1110101101:	sigmoid = 7'b0101100;
		10'b1110101110:	sigmoid = 7'b0101100;
		10'b1110101111:	sigmoid = 7'b0101100;
		10'b1110110000:	sigmoid = 7'b0101101;
		10'b1110110001:	sigmoid = 7'b0101101;
		10'b1110110010:	sigmoid = 7'b0101101;
		10'b1110110011:	sigmoid = 7'b0101101;
		10'b1110110100:	sigmoid = 7'b0101110;
		10'b1110110101:	sigmoid = 7'b0101110;
		10'b1110110110:	sigmoid = 7'b0101110;
		10'b1110110111:	sigmoid = 7'b0101110;
		10'b1110111000:	sigmoid = 7'b0101110;
		10'b1110111001:	sigmoid = 7'b0101111;
		10'b1110111010:	sigmoid = 7'b0101111;
		10'b1110111011:	sigmoid = 7'b0101111;
		10'b1110111100:	sigmoid = 7'b0101111;
		10'b1110111101:	sigmoid = 7'b0110000;
		10'b1110111110:	sigmoid = 7'b0110000;
		10'b1110111111:	sigmoid = 7'b0110000;
		10'b1111000000:	sigmoid = 7'b0110000;
		10'b1111000001:	sigmoid = 7'b0110001;
		10'b1111000010:	sigmoid = 7'b0110001;
		10'b1111000011:	sigmoid = 7'b0110001;
		10'b1111000100:	sigmoid = 7'b0110001;
		10'b1111000101:	sigmoid = 7'b0110010;
		10'b1111000110:	sigmoid = 7'b0110010;
		10'b1111000111:	sigmoid = 7'b0110010;
		10'b1111001000:	sigmoid = 7'b0110010;
		10'b1111001001:	sigmoid = 7'b0110010;
		10'b1111001010:	sigmoid = 7'b0110011;
		10'b1111001011:	sigmoid = 7'b0110011;
		10'b1111001100:	sigmoid = 7'b0110011;
		10'b1111001101:	sigmoid = 7'b0110011;
		10'b1111001110:	sigmoid = 7'b0110100;
		10'b1111001111:	sigmoid = 7'b0110100;
		10'b1111010000:	sigmoid = 7'b0110100;
		10'b1111010001:	sigmoid = 7'b0110100;
		10'b1111010010:	sigmoid = 7'b0110101;
		10'b1111010011:	sigmoid = 7'b0110101;
		10'b1111010100:	sigmoid = 7'b0110101;
		10'b1111010101:	sigmoid = 7'b0110101;
		10'b1111010110:	sigmoid = 7'b0110110;
		10'b1111010111:	sigmoid = 7'b0110110;
		10'b1111011000:	sigmoid = 7'b0110110;
		10'b1111011001:	sigmoid = 7'b0110110;
		10'b1111011010:	sigmoid = 7'b0110111;
		10'b1111011011:	sigmoid = 7'b0110111;
		10'b1111011100:	sigmoid = 7'b0110111;
		10'b1111011101:	sigmoid = 7'b0110111;
		10'b1111011110:	sigmoid = 7'b0111000;
		10'b1111011111:	sigmoid = 7'b0111000;
		10'b1111100000:	sigmoid = 7'b0111000;
		10'b1111100001:	sigmoid = 7'b0111000;
		10'b1111100010:	sigmoid = 7'b0111001;
		10'b1111100011:	sigmoid = 7'b0111001;
		10'b1111100100:	sigmoid = 7'b0111001;
		10'b1111100101:	sigmoid = 7'b0111001;
		10'b1111100110:	sigmoid = 7'b0111010;
		10'b1111100111:	sigmoid = 7'b0111010;
		10'b1111101000:	sigmoid = 7'b0111010;
		10'b1111101001:	sigmoid = 7'b0111010;
		10'b1111101010:	sigmoid = 7'b0111011;
		10'b1111101011:	sigmoid = 7'b0111011;
		10'b1111101100:	sigmoid = 7'b0111011;
		10'b1111101101:	sigmoid = 7'b0111011;
		10'b1111101110:	sigmoid = 7'b0111100;
		10'b1111101111:	sigmoid = 7'b0111100;
		10'b1111110000:	sigmoid = 7'b0111100;
		10'b1111110001:	sigmoid = 7'b0111100;
		10'b1111110010:	sigmoid = 7'b0111101;
		10'b1111110011:	sigmoid = 7'b0111101;
		10'b1111110100:	sigmoid = 7'b0111101;
		10'b1111110101:	sigmoid = 7'b0111101;
		10'b1111110110:	sigmoid = 7'b0111110;
		10'b1111110111:	sigmoid = 7'b0111110;
		10'b1111111000:	sigmoid = 7'b0111110;
		10'b1111111001:	sigmoid = 7'b0111110;
		10'b1111111010:	sigmoid = 7'b0111111;
		10'b1111111011:	sigmoid = 7'b0111111;
		10'b1111111100:	sigmoid = 7'b0111111;
		10'b1111111101:	sigmoid = 7'b0111111;
		10'b1111111110:	sigmoid = 7'b1000000;
		10'b1111111111:	sigmoid = 7'b1000000;
		10'b0000000000:	sigmoid = 7'b1000000;
		10'b0000000001:	sigmoid = 7'b1000000;
		10'b0000000010:	sigmoid = 7'b1000000;
		10'b0000000011:	sigmoid = 7'b1000001;
		10'b0000000100:	sigmoid = 7'b1000001;
		10'b0000000101:	sigmoid = 7'b1000001;
		10'b0000000110:	sigmoid = 7'b1000001;
		10'b0000000111:	sigmoid = 7'b1000010;
		10'b0000001000:	sigmoid = 7'b1000010;
		10'b0000001001:	sigmoid = 7'b1000010;
		10'b0000001010:	sigmoid = 7'b1000010;
		10'b0000001011:	sigmoid = 7'b1000011;
		10'b0000001100:	sigmoid = 7'b1000011;
		10'b0000001101:	sigmoid = 7'b1000011;
		10'b0000001110:	sigmoid = 7'b1000011;
		10'b0000001111:	sigmoid = 7'b1000100;
		10'b0000010000:	sigmoid = 7'b1000100;
		10'b0000010001:	sigmoid = 7'b1000100;
		10'b0000010010:	sigmoid = 7'b1000100;
		10'b0000010011:	sigmoid = 7'b1000101;
		10'b0000010100:	sigmoid = 7'b1000101;
		10'b0000010101:	sigmoid = 7'b1000101;
		10'b0000010110:	sigmoid = 7'b1000101;
		10'b0000010111:	sigmoid = 7'b1000110;
		10'b0000011000:	sigmoid = 7'b1000110;
		10'b0000011001:	sigmoid = 7'b1000110;
		10'b0000011010:	sigmoid = 7'b1000110;
		10'b0000011011:	sigmoid = 7'b1000111;
		10'b0000011100:	sigmoid = 7'b1000111;
		10'b0000011101:	sigmoid = 7'b1000111;
		10'b0000011110:	sigmoid = 7'b1000111;
		10'b0000011111:	sigmoid = 7'b1001000;
		10'b0000100000:	sigmoid = 7'b1001000;
		10'b0000100001:	sigmoid = 7'b1001000;
		10'b0000100010:	sigmoid = 7'b1001000;
		10'b0000100011:	sigmoid = 7'b1001001;
		10'b0000100100:	sigmoid = 7'b1001001;
		10'b0000100101:	sigmoid = 7'b1001001;
		10'b0000100110:	sigmoid = 7'b1001001;
		10'b0000100111:	sigmoid = 7'b1001010;
		10'b0000101000:	sigmoid = 7'b1001010;
		10'b0000101001:	sigmoid = 7'b1001010;
		10'b0000101010:	sigmoid = 7'b1001010;
		10'b0000101011:	sigmoid = 7'b1001011;
		10'b0000101100:	sigmoid = 7'b1001011;
		10'b0000101101:	sigmoid = 7'b1001011;
		10'b0000101110:	sigmoid = 7'b1001011;
		10'b0000101111:	sigmoid = 7'b1001100;
		10'b0000110000:	sigmoid = 7'b1001100;
		10'b0000110001:	sigmoid = 7'b1001100;
		10'b0000110010:	sigmoid = 7'b1001100;
		10'b0000110011:	sigmoid = 7'b1001101;
		10'b0000110100:	sigmoid = 7'b1001101;
		10'b0000110101:	sigmoid = 7'b1001101;
		10'b0000110110:	sigmoid = 7'b1001101;
		10'b0000110111:	sigmoid = 7'b1001110;
		10'b0000111000:	sigmoid = 7'b1001110;
		10'b0000111001:	sigmoid = 7'b1001110;
		10'b0000111010:	sigmoid = 7'b1001110;
		10'b0000111011:	sigmoid = 7'b1001110;
		10'b0000111100:	sigmoid = 7'b1001111;
		10'b0000111101:	sigmoid = 7'b1001111;
		10'b0000111110:	sigmoid = 7'b1001111;
		10'b0000111111:	sigmoid = 7'b1001111;
		10'b0001000000:	sigmoid = 7'b1010000;
		10'b0001000001:	sigmoid = 7'b1010000;
		10'b0001000010:	sigmoid = 7'b1010000;
		10'b0001000011:	sigmoid = 7'b1010000;
		10'b0001000100:	sigmoid = 7'b1010001;
		10'b0001000101:	sigmoid = 7'b1010001;
		10'b0001000110:	sigmoid = 7'b1010001;
		10'b0001000111:	sigmoid = 7'b1010001;
		10'b0001001000:	sigmoid = 7'b1010010;
		10'b0001001001:	sigmoid = 7'b1010010;
		10'b0001001010:	sigmoid = 7'b1010010;
		10'b0001001011:	sigmoid = 7'b1010010;
		10'b0001001100:	sigmoid = 7'b1010010;
		10'b0001001101:	sigmoid = 7'b1010011;
		10'b0001001110:	sigmoid = 7'b1010011;
		10'b0001001111:	sigmoid = 7'b1010011;
		10'b0001010000:	sigmoid = 7'b1010011;
		10'b0001010001:	sigmoid = 7'b1010100;
		10'b0001010010:	sigmoid = 7'b1010100;
		10'b0001010011:	sigmoid = 7'b1010100;
		10'b0001010100:	sigmoid = 7'b1010100;
		10'b0001010101:	sigmoid = 7'b1010101;
		10'b0001010110:	sigmoid = 7'b1010101;
		10'b0001010111:	sigmoid = 7'b1010101;
		10'b0001011000:	sigmoid = 7'b1010101;
		10'b0001011001:	sigmoid = 7'b1010101;
		10'b0001011010:	sigmoid = 7'b1010110;
		10'b0001011011:	sigmoid = 7'b1010110;
		10'b0001011100:	sigmoid = 7'b1010110;
		10'b0001011101:	sigmoid = 7'b1010110;
		10'b0001011110:	sigmoid = 7'b1010110;
		10'b0001011111:	sigmoid = 7'b1010111;
		10'b0001100000:	sigmoid = 7'b1010111;
		10'b0001100001:	sigmoid = 7'b1010111;
		10'b0001100010:	sigmoid = 7'b1010111;
		10'b0001100011:	sigmoid = 7'b1011000;
		10'b0001100100:	sigmoid = 7'b1011000;
		10'b0001100101:	sigmoid = 7'b1011000;
		10'b0001100110:	sigmoid = 7'b1011000;
		10'b0001100111:	sigmoid = 7'b1011000;
		10'b0001101000:	sigmoid = 7'b1011001;
		10'b0001101001:	sigmoid = 7'b1011001;
		10'b0001101010:	sigmoid = 7'b1011001;
		10'b0001101011:	sigmoid = 7'b1011001;
		10'b0001101100:	sigmoid = 7'b1011010;
		10'b0001101101:	sigmoid = 7'b1011010;
		10'b0001101110:	sigmoid = 7'b1011010;
		10'b0001101111:	sigmoid = 7'b1011010;
		10'b0001110000:	sigmoid = 7'b1011010;
		10'b0001110001:	sigmoid = 7'b1011011;
		10'b0001110010:	sigmoid = 7'b1011011;
		10'b0001110011:	sigmoid = 7'b1011011;
		10'b0001110100:	sigmoid = 7'b1011011;
		10'b0001110101:	sigmoid = 7'b1011011;
		10'b0001110110:	sigmoid = 7'b1011100;
		10'b0001110111:	sigmoid = 7'b1011100;
		10'b0001111000:	sigmoid = 7'b1011100;
		10'b0001111001:	sigmoid = 7'b1011100;
		10'b0001111010:	sigmoid = 7'b1011100;
		10'b0001111011:	sigmoid = 7'b1011101;
		10'b0001111100:	sigmoid = 7'b1011101;
		10'b0001111101:	sigmoid = 7'b1011101;
		10'b0001111110:	sigmoid = 7'b1011101;
		10'b0001111111:	sigmoid = 7'b1011101;
		10'b0010000000:	sigmoid = 7'b1011110;
		10'b0010000001:	sigmoid = 7'b1011110;
		10'b0010000010:	sigmoid = 7'b1011110;
		10'b0010000011:	sigmoid = 7'b1011110;
		10'b0010000100:	sigmoid = 7'b1011110;
		10'b0010000101:	sigmoid = 7'b1011111;
		10'b0010000110:	sigmoid = 7'b1011111;
		10'b0010000111:	sigmoid = 7'b1011111;
		10'b0010001000:	sigmoid = 7'b1011111;
		10'b0010001001:	sigmoid = 7'b1011111;
		10'b0010001010:	sigmoid = 7'b1100000;
		10'b0010001011:	sigmoid = 7'b1100000;
		10'b0010001100:	sigmoid = 7'b1100000;
		10'b0010001101:	sigmoid = 7'b1100000;
		10'b0010001110:	sigmoid = 7'b1100000;
		10'b0010001111:	sigmoid = 7'b1100000;
		10'b0010010000:	sigmoid = 7'b1100001;
		10'b0010010001:	sigmoid = 7'b1100001;
		10'b0010010010:	sigmoid = 7'b1100001;
		10'b0010010011:	sigmoid = 7'b1100001;
		10'b0010010100:	sigmoid = 7'b1100001;
		10'b0010010101:	sigmoid = 7'b1100010;
		10'b0010010110:	sigmoid = 7'b1100010;
		10'b0010010111:	sigmoid = 7'b1100010;
		10'b0010011000:	sigmoid = 7'b1100010;
		10'b0010011001:	sigmoid = 7'b1100010;
		10'b0010011010:	sigmoid = 7'b1100010;
		10'b0010011011:	sigmoid = 7'b1100011;
		10'b0010011100:	sigmoid = 7'b1100011;
		10'b0010011101:	sigmoid = 7'b1100011;
		10'b0010011110:	sigmoid = 7'b1100011;
		10'b0010011111:	sigmoid = 7'b1100011;
		10'b0010100000:	sigmoid = 7'b1100011;
		10'b0010100001:	sigmoid = 7'b1100100;
		10'b0010100010:	sigmoid = 7'b1100100;
		10'b0010100011:	sigmoid = 7'b1100100;
		10'b0010100100:	sigmoid = 7'b1100100;
		10'b0010100101:	sigmoid = 7'b1100100;
		10'b0010100110:	sigmoid = 7'b1100101;
		10'b0010100111:	sigmoid = 7'b1100101;
		10'b0010101000:	sigmoid = 7'b1100101;
		10'b0010101001:	sigmoid = 7'b1100101;
		10'b0010101010:	sigmoid = 7'b1100101;
		10'b0010101011:	sigmoid = 7'b1100101;
		10'b0010101100:	sigmoid = 7'b1100110;
		10'b0010101101:	sigmoid = 7'b1100110;
		10'b0010101110:	sigmoid = 7'b1100110;
		10'b0010101111:	sigmoid = 7'b1100110;
		10'b0010110000:	sigmoid = 7'b1100110;
		10'b0010110001:	sigmoid = 7'b1100110;
		10'b0010110010:	sigmoid = 7'b1100110;
		10'b0010110011:	sigmoid = 7'b1100111;
		10'b0010110100:	sigmoid = 7'b1100111;
		10'b0010110101:	sigmoid = 7'b1100111;
		10'b0010110110:	sigmoid = 7'b1100111;
		10'b0010110111:	sigmoid = 7'b1100111;
		10'b0010111000:	sigmoid = 7'b1100111;
		10'b0010111001:	sigmoid = 7'b1101000;
		10'b0010111010:	sigmoid = 7'b1101000;
		10'b0010111011:	sigmoid = 7'b1101000;
		10'b0010111100:	sigmoid = 7'b1101000;
		10'b0010111101:	sigmoid = 7'b1101000;
		10'b0010111110:	sigmoid = 7'b1101000;
		10'b0010111111:	sigmoid = 7'b1101001;
		10'b0011000000:	sigmoid = 7'b1101001;
		10'b0011000001:	sigmoid = 7'b1101001;
		10'b0011000010:	sigmoid = 7'b1101001;
		10'b0011000011:	sigmoid = 7'b1101001;
		10'b0011000100:	sigmoid = 7'b1101001;
		10'b0011000101:	sigmoid = 7'b1101001;
		10'b0011000110:	sigmoid = 7'b1101010;
		10'b0011000111:	sigmoid = 7'b1101010;
		10'b0011001000:	sigmoid = 7'b1101010;
		10'b0011001001:	sigmoid = 7'b1101010;
		10'b0011001010:	sigmoid = 7'b1101010;
		10'b0011001011:	sigmoid = 7'b1101010;
		10'b0011001100:	sigmoid = 7'b1101010;
		10'b0011001101:	sigmoid = 7'b1101011;
		10'b0011001110:	sigmoid = 7'b1101011;
		10'b0011001111:	sigmoid = 7'b1101011;
		10'b0011010000:	sigmoid = 7'b1101011;
		10'b0011010001:	sigmoid = 7'b1101011;
		10'b0011010010:	sigmoid = 7'b1101011;
		10'b0011010011:	sigmoid = 7'b1101011;
		10'b0011010100:	sigmoid = 7'b1101011;
		10'b0011010101:	sigmoid = 7'b1101100;
		10'b0011010110:	sigmoid = 7'b1101100;
		10'b0011010111:	sigmoid = 7'b1101100;
		10'b0011011000:	sigmoid = 7'b1101100;
		10'b0011011001:	sigmoid = 7'b1101100;
		10'b0011011010:	sigmoid = 7'b1101100;
		10'b0011011011:	sigmoid = 7'b1101100;
		10'b0011011100:	sigmoid = 7'b1101101;
		10'b0011011101:	sigmoid = 7'b1101101;
		10'b0011011110:	sigmoid = 7'b1101101;
		10'b0011011111:	sigmoid = 7'b1101101;
		10'b0011100000:	sigmoid = 7'b1101101;
		10'b0011100001:	sigmoid = 7'b1101101;
		10'b0011100010:	sigmoid = 7'b1101101;
		10'b0011100011:	sigmoid = 7'b1101101;
		10'b0011100100:	sigmoid = 7'b1101110;
		10'b0011100101:	sigmoid = 7'b1101110;
		10'b0011100110:	sigmoid = 7'b1101110;
		10'b0011100111:	sigmoid = 7'b1101110;
		10'b0011101000:	sigmoid = 7'b1101110;
		10'b0011101001:	sigmoid = 7'b1101110;
		10'b0011101010:	sigmoid = 7'b1101110;
		10'b0011101011:	sigmoid = 7'b1101110;
		10'b0011101100:	sigmoid = 7'b1101111;
		10'b0011101101:	sigmoid = 7'b1101111;
		10'b0011101110:	sigmoid = 7'b1101111;
		10'b0011101111:	sigmoid = 7'b1101111;
		10'b0011110000:	sigmoid = 7'b1101111;
		10'b0011110001:	sigmoid = 7'b1101111;
		10'b0011110010:	sigmoid = 7'b1101111;
		10'b0011110011:	sigmoid = 7'b1101111;
		10'b0011110100:	sigmoid = 7'b1101111;
		10'b0011110101:	sigmoid = 7'b1110000;
		10'b0011110110:	sigmoid = 7'b1110000;
		10'b0011110111:	sigmoid = 7'b1110000;
		10'b0011111000:	sigmoid = 7'b1110000;
		10'b0011111001:	sigmoid = 7'b1110000;
		10'b0011111010:	sigmoid = 7'b1110000;
		10'b0011111011:	sigmoid = 7'b1110000;
		10'b0011111100:	sigmoid = 7'b1110000;
		10'b0011111101:	sigmoid = 7'b1110000;
		10'b0011111110:	sigmoid = 7'b1110001;
		10'b0011111111:	sigmoid = 7'b1110001;
		10'b0100000000:	sigmoid = 7'b1110001;
		10'b0100000001:	sigmoid = 7'b1110001;
		10'b0100000010:	sigmoid = 7'b1110001;
		10'b0100000011:	sigmoid = 7'b1110001;
		10'b0100000100:	sigmoid = 7'b1110001;
		10'b0100000101:	sigmoid = 7'b1110001;
		10'b0100000110:	sigmoid = 7'b1110001;
		10'b0100000111:	sigmoid = 7'b1110001;
		10'b0100001000:	sigmoid = 7'b1110010;
		10'b0100001001:	sigmoid = 7'b1110010;
		10'b0100001010:	sigmoid = 7'b1110010;
		10'b0100001011:	sigmoid = 7'b1110010;
		10'b0100001100:	sigmoid = 7'b1110010;
		10'b0100001101:	sigmoid = 7'b1110010;
		10'b0100001110:	sigmoid = 7'b1110010;
		10'b0100001111:	sigmoid = 7'b1110010;
		10'b0100010000:	sigmoid = 7'b1110010;
		10'b0100010001:	sigmoid = 7'b1110010;
		10'b0100010010:	sigmoid = 7'b1110011;
		10'b0100010011:	sigmoid = 7'b1110011;
		10'b0100010100:	sigmoid = 7'b1110011;
		10'b0100010101:	sigmoid = 7'b1110011;
		10'b0100010110:	sigmoid = 7'b1110011;
		10'b0100010111:	sigmoid = 7'b1110011;
		10'b0100011000:	sigmoid = 7'b1110011;
		10'b0100011001:	sigmoid = 7'b1110011;
		10'b0100011010:	sigmoid = 7'b1110011;
		10'b0100011011:	sigmoid = 7'b1110011;
		10'b0100011100:	sigmoid = 7'b1110011;
		10'b0100011101:	sigmoid = 7'b1110100;
		10'b0100011110:	sigmoid = 7'b1110100;
		10'b0100011111:	sigmoid = 7'b1110100;
		10'b0100100000:	sigmoid = 7'b1110100;
		10'b0100100001:	sigmoid = 7'b1110100;
		10'b0100100010:	sigmoid = 7'b1110100;
		10'b0100100011:	sigmoid = 7'b1110100;
		10'b0100100100:	sigmoid = 7'b1110100;
		10'b0100100101:	sigmoid = 7'b1110100;
		10'b0100100110:	sigmoid = 7'b1110100;
		10'b0100100111:	sigmoid = 7'b1110100;
		10'b0100101000:	sigmoid = 7'b1110100;
		10'b0100101001:	sigmoid = 7'b1110101;
		10'b0100101010:	sigmoid = 7'b1110101;
		10'b0100101011:	sigmoid = 7'b1110101;
		10'b0100101100:	sigmoid = 7'b1110101;
		10'b0100101101:	sigmoid = 7'b1110101;
		10'b0100101110:	sigmoid = 7'b1110101;
		10'b0100101111:	sigmoid = 7'b1110101;
		10'b0100110000:	sigmoid = 7'b1110101;
		10'b0100110001:	sigmoid = 7'b1110101;
		10'b0100110010:	sigmoid = 7'b1110101;
		10'b0100110011:	sigmoid = 7'b1110101;
		10'b0100110100:	sigmoid = 7'b1110101;
		10'b0100110101:	sigmoid = 7'b1110101;
		10'b0100110110:	sigmoid = 7'b1110110;
		10'b0100110111:	sigmoid = 7'b1110110;
		10'b0100111000:	sigmoid = 7'b1110110;
		10'b0100111001:	sigmoid = 7'b1110110;
		10'b0100111010:	sigmoid = 7'b1110110;
		10'b0100111011:	sigmoid = 7'b1110110;
		10'b0100111100:	sigmoid = 7'b1110110;
		10'b0100111101:	sigmoid = 7'b1110110;
		10'b0100111110:	sigmoid = 7'b1110110;
		10'b0100111111:	sigmoid = 7'b1110110;
		10'b0101000000:	sigmoid = 7'b1110110;
		10'b0101000001:	sigmoid = 7'b1110110;
		10'b0101000010:	sigmoid = 7'b1110110;
		10'b0101000011:	sigmoid = 7'b1110110;
		10'b0101000100:	sigmoid = 7'b1110111;
		10'b0101000101:	sigmoid = 7'b1110111;
		10'b0101000110:	sigmoid = 7'b1110111;
		10'b0101000111:	sigmoid = 7'b1110111;
		10'b0101001000:	sigmoid = 7'b1110111;
		10'b0101001001:	sigmoid = 7'b1110111;
		10'b0101001010:	sigmoid = 7'b1110111;
		10'b0101001011:	sigmoid = 7'b1110111;
		10'b0101001100:	sigmoid = 7'b1110111;
		10'b0101001101:	sigmoid = 7'b1110111;
		10'b0101001110:	sigmoid = 7'b1110111;
		10'b0101001111:	sigmoid = 7'b1110111;
		10'b0101010000:	sigmoid = 7'b1110111;
		10'b0101010001:	sigmoid = 7'b1110111;
		10'b0101010010:	sigmoid = 7'b1110111;
		10'b0101010011:	sigmoid = 7'b1111000;
		10'b0101010100:	sigmoid = 7'b1111000;
		10'b0101010101:	sigmoid = 7'b1111000;
		10'b0101010110:	sigmoid = 7'b1111000;
		10'b0101010111:	sigmoid = 7'b1111000;
		10'b0101011000:	sigmoid = 7'b1111000;
		10'b0101011001:	sigmoid = 7'b1111000;
		10'b0101011010:	sigmoid = 7'b1111000;
		10'b0101011011:	sigmoid = 7'b1111000;
		10'b0101011100:	sigmoid = 7'b1111000;
		10'b0101011101:	sigmoid = 7'b1111000;
		10'b0101011110:	sigmoid = 7'b1111000;
		10'b0101011111:	sigmoid = 7'b1111000;
		10'b0101100000:	sigmoid = 7'b1111000;
		10'b0101100001:	sigmoid = 7'b1111000;
		10'b0101100010:	sigmoid = 7'b1111000;
		10'b0101100011:	sigmoid = 7'b1111000;
		10'b0101100100:	sigmoid = 7'b1111001;
		10'b0101100101:	sigmoid = 7'b1111001;
		10'b0101100110:	sigmoid = 7'b1111001;
		10'b0101100111:	sigmoid = 7'b1111001;
		10'b0101101000:	sigmoid = 7'b1111001;
		10'b0101101001:	sigmoid = 7'b1111001;
		10'b0101101010:	sigmoid = 7'b1111001;
		10'b0101101011:	sigmoid = 7'b1111001;
		10'b0101101100:	sigmoid = 7'b1111001;
		10'b0101101101:	sigmoid = 7'b1111001;
		10'b0101101110:	sigmoid = 7'b1111001;
		10'b0101101111:	sigmoid = 7'b1111001;
		10'b0101110000:	sigmoid = 7'b1111001;
		10'b0101110001:	sigmoid = 7'b1111001;
		10'b0101110010:	sigmoid = 7'b1111001;
		10'b0101110011:	sigmoid = 7'b1111001;
		10'b0101110100:	sigmoid = 7'b1111001;
		10'b0101110101:	sigmoid = 7'b1111001;
		10'b0101110110:	sigmoid = 7'b1111001;
		10'b0101110111:	sigmoid = 7'b1111010;
		10'b0101111000:	sigmoid = 7'b1111010;
		10'b0101111001:	sigmoid = 7'b1111010;
		10'b0101111010:	sigmoid = 7'b1111010;
		10'b0101111011:	sigmoid = 7'b1111010;
		10'b0101111100:	sigmoid = 7'b1111010;
		10'b0101111101:	sigmoid = 7'b1111010;
		10'b0101111110:	sigmoid = 7'b1111010;
		10'b0101111111:	sigmoid = 7'b1111010;
		10'b0110000000:	sigmoid = 7'b1111010;
		10'b0110000001:	sigmoid = 7'b1111010;
		10'b0110000010:	sigmoid = 7'b1111010;
		10'b0110000011:	sigmoid = 7'b1111010;
		10'b0110000100:	sigmoid = 7'b1111010;
		10'b0110000101:	sigmoid = 7'b1111010;
		10'b0110000110:	sigmoid = 7'b1111010;
		10'b0110000111:	sigmoid = 7'b1111010;
		10'b0110001000:	sigmoid = 7'b1111010;
		10'b0110001001:	sigmoid = 7'b1111010;
		10'b0110001010:	sigmoid = 7'b1111010;
		10'b0110001011:	sigmoid = 7'b1111010;
		10'b0110001100:	sigmoid = 7'b1111010;
		10'b0110001101:	sigmoid = 7'b1111010;
		10'b0110001110:	sigmoid = 7'b1111011;
		10'b0110001111:	sigmoid = 7'b1111011;
		10'b0110010000:	sigmoid = 7'b1111011;
		10'b0110010001:	sigmoid = 7'b1111011;
		10'b0110010010:	sigmoid = 7'b1111011;
		10'b0110010011:	sigmoid = 7'b1111011;
		10'b0110010100:	sigmoid = 7'b1111011;
		10'b0110010101:	sigmoid = 7'b1111011;
		10'b0110010110:	sigmoid = 7'b1111011;
		10'b0110010111:	sigmoid = 7'b1111011;
		10'b0110011000:	sigmoid = 7'b1111011;
		10'b0110011001:	sigmoid = 7'b1111011;
		10'b0110011010:	sigmoid = 7'b1111011;
		10'b0110011011:	sigmoid = 7'b1111011;
		10'b0110011100:	sigmoid = 7'b1111011;
		10'b0110011101:	sigmoid = 7'b1111011;
		10'b0110011110:	sigmoid = 7'b1111011;
		10'b0110011111:	sigmoid = 7'b1111011;
		10'b0110100000:	sigmoid = 7'b1111011;
		10'b0110100001:	sigmoid = 7'b1111011;
		10'b0110100010:	sigmoid = 7'b1111011;
		10'b0110100011:	sigmoid = 7'b1111011;
		10'b0110100100:	sigmoid = 7'b1111011;
		10'b0110100101:	sigmoid = 7'b1111011;
		10'b0110100110:	sigmoid = 7'b1111011;
		10'b0110100111:	sigmoid = 7'b1111011;
		10'b0110101000:	sigmoid = 7'b1111100;
		10'b0110101001:	sigmoid = 7'b1111100;
		10'b0110101010:	sigmoid = 7'b1111100;
		10'b0110101011:	sigmoid = 7'b1111100;
		10'b0110101100:	sigmoid = 7'b1111100;
		10'b0110101101:	sigmoid = 7'b1111100;
		10'b0110101110:	sigmoid = 7'b1111100;
		10'b0110101111:	sigmoid = 7'b1111100;
		10'b0110110000:	sigmoid = 7'b1111100;
		10'b0110110001:	sigmoid = 7'b1111100;
		10'b0110110010:	sigmoid = 7'b1111100;
		10'b0110110011:	sigmoid = 7'b1111100;
		10'b0110110100:	sigmoid = 7'b1111100;
		10'b0110110101:	sigmoid = 7'b1111100;
		10'b0110110110:	sigmoid = 7'b1111100;
		10'b0110110111:	sigmoid = 7'b1111100;
		10'b0110111000:	sigmoid = 7'b1111100;
		10'b0110111001:	sigmoid = 7'b1111100;
		10'b0110111010:	sigmoid = 7'b1111100;
		10'b0110111011:	sigmoid = 7'b1111100;
		10'b0110111100:	sigmoid = 7'b1111100;
		10'b0110111101:	sigmoid = 7'b1111100;
		10'b0110111110:	sigmoid = 7'b1111100;
		10'b0110111111:	sigmoid = 7'b1111100;
		10'b0111000000:	sigmoid = 7'b1111100;
		10'b0111000001:	sigmoid = 7'b1111100;
		10'b0111000010:	sigmoid = 7'b1111100;
		10'b0111000011:	sigmoid = 7'b1111100;
		10'b0111000100:	sigmoid = 7'b1111100;
		10'b0111000101:	sigmoid = 7'b1111100;
		10'b0111000110:	sigmoid = 7'b1111100;
		10'b0111000111:	sigmoid = 7'b1111100;
		10'b0111001000:	sigmoid = 7'b1111100;
		10'b0111001001:	sigmoid = 7'b1111100;
		10'b0111001010:	sigmoid = 7'b1111101;
		10'b0111001011:	sigmoid = 7'b1111101;
		10'b0111001100:	sigmoid = 7'b1111101;
		10'b0111001101:	sigmoid = 7'b1111101;
		10'b0111001110:	sigmoid = 7'b1111101;
		10'b0111001111:	sigmoid = 7'b1111101;
		10'b0111010000:	sigmoid = 7'b1111101;
		10'b0111010001:	sigmoid = 7'b1111101;
		10'b0111010010:	sigmoid = 7'b1111101;
		10'b0111010011:	sigmoid = 7'b1111101;
		10'b0111010100:	sigmoid = 7'b1111101;
		10'b0111010101:	sigmoid = 7'b1111101;
		10'b0111010110:	sigmoid = 7'b1111101;
		10'b0111010111:	sigmoid = 7'b1111101;
		10'b0111011000:	sigmoid = 7'b1111101;
		10'b0111011001:	sigmoid = 7'b1111101;
		10'b0111011010:	sigmoid = 7'b1111101;
		10'b0111011011:	sigmoid = 7'b1111101;
		10'b0111011100:	sigmoid = 7'b1111101;
		10'b0111011101:	sigmoid = 7'b1111101;
		10'b0111011110:	sigmoid = 7'b1111101;
		10'b0111011111:	sigmoid = 7'b1111101;
		10'b0111100000:	sigmoid = 7'b1111101;
		10'b0111100001:	sigmoid = 7'b1111101;
		10'b0111100010:	sigmoid = 7'b1111101;
		10'b0111100011:	sigmoid = 7'b1111101;
		10'b0111100100:	sigmoid = 7'b1111101;
		10'b0111100101:	sigmoid = 7'b1111101;
		10'b0111100110:	sigmoid = 7'b1111101;
		10'b0111100111:	sigmoid = 7'b1111101;
		10'b0111101000:	sigmoid = 7'b1111101;
		10'b0111101001:	sigmoid = 7'b1111101;
		10'b0111101010:	sigmoid = 7'b1111101;
		10'b0111101011:	sigmoid = 7'b1111101;
		10'b0111101100:	sigmoid = 7'b1111101;
		10'b0111101101:	sigmoid = 7'b1111101;
		10'b0111101110:	sigmoid = 7'b1111101;
		10'b0111101111:	sigmoid = 7'b1111101;
		10'b0111110000:	sigmoid = 7'b1111101;
		10'b0111110001:	sigmoid = 7'b1111101;
		10'b0111110010:	sigmoid = 7'b1111101;
		10'b0111110011:	sigmoid = 7'b1111101;
		10'b0111110100:	sigmoid = 7'b1111101;
		10'b0111110101:	sigmoid = 7'b1111101;
		10'b0111110110:	sigmoid = 7'b1111110;
		10'b0111110111:	sigmoid = 7'b1111110;
		10'b0111111000:	sigmoid = 7'b1111110;
		10'b0111111001:	sigmoid = 7'b1111110;
		10'b0111111010:	sigmoid = 7'b1111110;
		10'b0111111011:	sigmoid = 7'b1111110;
		10'b0111111100:	sigmoid = 7'b1111110;
		10'b0111111101:	sigmoid = 7'b1111110;
		10'b0111111110:	sigmoid = 7'b1111110;
		10'b0111111111:	sigmoid = 7'b1111110;

	endcase
endmodule

// __________________________________________________________________________________________________________ //
// __________________________________________________________________________________________________________ //

module sig_prime #(
	parameter width = 10, 
	parameter int_bits = 2,
	parameter frac_bits = width-int_bits-1,
	parameter maxdomain = (2**int_bits>8) ? 8 : 2**int_bits,
	parameter lut_size = (2**width>4096) ? 4096 : 2**width
)(
	input clk,
	input signed [width-1:0] z,
	output reg[width-1:0] sp_out
);

	reg [frac_bits-3:0] sigmoid_prime; //since 2 MSB in frac_part are always 00

	/*always @(posedge clk)
	if(z[width-1]==1||z==0)
		sp_out = (z[width-1:width-int_bits+2] == 0 ||&z[width-1:width-int_bits+2])? 
			{{(int_bits+1){1'b0}},sigmoid_prime,3'b0}:1;//0;
	else
		//sp_out = (z[width-1:width-int_bits+2] == 0 ||&z[width-1:width-int_bits+2])? 
		//	{{(int_bits+1){1'b0}},sigmoid_prime,3'b0}:1;
		sp_out = 1'b1<<frac_bits;*/
	
	
	always @(posedge clk) begin
		sp_out = (z[width-1:width-int_bits+$clog2(maxdomain)-1] == 0 || &z[width-1:width-int_bits+$clog2(maxdomain)-1]) ? 
		{{(int_bits+3){1'b0}},sigmoid_prime} : //since 2 MSB in frac_part are always 00
		1; //If z is outside [-maxdomain,+maxdomain], sigmoid prime will always be 0. This is stored as all zeros followed by 1 at LSB, i.e. 2^(-frac_bits), which is the lowest number possible (~=0)
	end

	always @(z[frac_bits+$clog2(maxdomain):frac_bits-$clog2(lut_size)+$clog2(maxdomain)+1]) //this ensures that we read exactly log(lut_size) bits as address of LUT
	case (z[frac_bits+$clog2(maxdomain):frac_bits-$clog2(lut_size)+$clog2(maxdomain)+1])
		
		10'b1000000000:	sigmoid_prime = 5'b00010;
		10'b1000000001:	sigmoid_prime = 5'b00010;
		10'b1000000010:	sigmoid_prime = 5'b00010;
		10'b1000000011:	sigmoid_prime = 5'b00010;
		10'b1000000100:	sigmoid_prime = 5'b00010;
		10'b1000000101:	sigmoid_prime = 5'b00010;
		10'b1000000110:	sigmoid_prime = 5'b00010;
		10'b1000000111:	sigmoid_prime = 5'b00010;
		10'b1000001000:	sigmoid_prime = 5'b00010;
		10'b1000001001:	sigmoid_prime = 5'b00010;
		10'b1000001010:	sigmoid_prime = 5'b00010;
		10'b1000001011:	sigmoid_prime = 5'b00010;
		10'b1000001100:	sigmoid_prime = 5'b00010;
		10'b1000001101:	sigmoid_prime = 5'b00010;
		10'b1000001110:	sigmoid_prime = 5'b00011;
		10'b1000001111:	sigmoid_prime = 5'b00011;
		10'b1000010000:	sigmoid_prime = 5'b00011;
		10'b1000010001:	sigmoid_prime = 5'b00011;
		10'b1000010010:	sigmoid_prime = 5'b00011;
		10'b1000010011:	sigmoid_prime = 5'b00011;
		10'b1000010100:	sigmoid_prime = 5'b00011;
		10'b1000010101:	sigmoid_prime = 5'b00011;
		10'b1000010110:	sigmoid_prime = 5'b00011;
		10'b1000010111:	sigmoid_prime = 5'b00011;
		10'b1000011000:	sigmoid_prime = 5'b00011;
		10'b1000011001:	sigmoid_prime = 5'b00011;
		10'b1000011010:	sigmoid_prime = 5'b00011;
		10'b1000011011:	sigmoid_prime = 5'b00011;
		10'b1000011100:	sigmoid_prime = 5'b00011;
		10'b1000011101:	sigmoid_prime = 5'b00011;
		10'b1000011110:	sigmoid_prime = 5'b00011;
		10'b1000011111:	sigmoid_prime = 5'b00011;
		10'b1000100000:	sigmoid_prime = 5'b00011;
		10'b1000100001:	sigmoid_prime = 5'b00011;
		10'b1000100010:	sigmoid_prime = 5'b00011;
		10'b1000100011:	sigmoid_prime = 5'b00011;
		10'b1000100100:	sigmoid_prime = 5'b00011;
		10'b1000100101:	sigmoid_prime = 5'b00011;
		10'b1000100110:	sigmoid_prime = 5'b00011;
		10'b1000100111:	sigmoid_prime = 5'b00011;
		10'b1000101000:	sigmoid_prime = 5'b00011;
		10'b1000101001:	sigmoid_prime = 5'b00011;
		10'b1000101010:	sigmoid_prime = 5'b00011;
		10'b1000101011:	sigmoid_prime = 5'b00011;
		10'b1000101100:	sigmoid_prime = 5'b00011;
		10'b1000101101:	sigmoid_prime = 5'b00011;
		10'b1000101110:	sigmoid_prime = 5'b00011;
		10'b1000101111:	sigmoid_prime = 5'b00011;
		10'b1000110000:	sigmoid_prime = 5'b00011;
		10'b1000110001:	sigmoid_prime = 5'b00011;
		10'b1000110010:	sigmoid_prime = 5'b00011;
		10'b1000110011:	sigmoid_prime = 5'b00011;
		10'b1000110100:	sigmoid_prime = 5'b00011;
		10'b1000110101:	sigmoid_prime = 5'b00011;
		10'b1000110110:	sigmoid_prime = 5'b00011;
		10'b1000110111:	sigmoid_prime = 5'b00011;
		10'b1000111000:	sigmoid_prime = 5'b00011;
		10'b1000111001:	sigmoid_prime = 5'b00011;
		10'b1000111010:	sigmoid_prime = 5'b00011;
		10'b1000111011:	sigmoid_prime = 5'b00100;
		10'b1000111100:	sigmoid_prime = 5'b00100;
		10'b1000111101:	sigmoid_prime = 5'b00100;
		10'b1000111110:	sigmoid_prime = 5'b00100;
		10'b1000111111:	sigmoid_prime = 5'b00100;
		10'b1001000000:	sigmoid_prime = 5'b00100;
		10'b1001000001:	sigmoid_prime = 5'b00100;
		10'b1001000010:	sigmoid_prime = 5'b00100;
		10'b1001000011:	sigmoid_prime = 5'b00100;
		10'b1001000100:	sigmoid_prime = 5'b00100;
		10'b1001000101:	sigmoid_prime = 5'b00100;
		10'b1001000110:	sigmoid_prime = 5'b00100;
		10'b1001000111:	sigmoid_prime = 5'b00100;
		10'b1001001000:	sigmoid_prime = 5'b00100;
		10'b1001001001:	sigmoid_prime = 5'b00100;
		10'b1001001010:	sigmoid_prime = 5'b00100;
		10'b1001001011:	sigmoid_prime = 5'b00100;
		10'b1001001100:	sigmoid_prime = 5'b00100;
		10'b1001001101:	sigmoid_prime = 5'b00100;
		10'b1001001110:	sigmoid_prime = 5'b00100;
		10'b1001001111:	sigmoid_prime = 5'b00100;
		10'b1001010000:	sigmoid_prime = 5'b00100;
		10'b1001010001:	sigmoid_prime = 5'b00100;
		10'b1001010010:	sigmoid_prime = 5'b00100;
		10'b1001010011:	sigmoid_prime = 5'b00100;
		10'b1001010100:	sigmoid_prime = 5'b00100;
		10'b1001010101:	sigmoid_prime = 5'b00100;
		10'b1001010110:	sigmoid_prime = 5'b00100;
		10'b1001010111:	sigmoid_prime = 5'b00100;
		10'b1001011000:	sigmoid_prime = 5'b00100;
		10'b1001011001:	sigmoid_prime = 5'b00100;
		10'b1001011010:	sigmoid_prime = 5'b00100;
		10'b1001011011:	sigmoid_prime = 5'b00100;
		10'b1001011100:	sigmoid_prime = 5'b00100;
		10'b1001011101:	sigmoid_prime = 5'b00101;
		10'b1001011110:	sigmoid_prime = 5'b00101;
		10'b1001011111:	sigmoid_prime = 5'b00101;
		10'b1001100000:	sigmoid_prime = 5'b00101;
		10'b1001100001:	sigmoid_prime = 5'b00101;
		10'b1001100010:	sigmoid_prime = 5'b00101;
		10'b1001100011:	sigmoid_prime = 5'b00101;
		10'b1001100100:	sigmoid_prime = 5'b00101;
		10'b1001100101:	sigmoid_prime = 5'b00101;
		10'b1001100110:	sigmoid_prime = 5'b00101;
		10'b1001100111:	sigmoid_prime = 5'b00101;
		10'b1001101000:	sigmoid_prime = 5'b00101;
		10'b1001101001:	sigmoid_prime = 5'b00101;
		10'b1001101010:	sigmoid_prime = 5'b00101;
		10'b1001101011:	sigmoid_prime = 5'b00101;
		10'b1001101100:	sigmoid_prime = 5'b00101;
		10'b1001101101:	sigmoid_prime = 5'b00101;
		10'b1001101110:	sigmoid_prime = 5'b00101;
		10'b1001101111:	sigmoid_prime = 5'b00101;
		10'b1001110000:	sigmoid_prime = 5'b00101;
		10'b1001110001:	sigmoid_prime = 5'b00101;
		10'b1001110010:	sigmoid_prime = 5'b00101;
		10'b1001110011:	sigmoid_prime = 5'b00101;
		10'b1001110100:	sigmoid_prime = 5'b00101;
		10'b1001110101:	sigmoid_prime = 5'b00101;
		10'b1001110110:	sigmoid_prime = 5'b00101;
		10'b1001110111:	sigmoid_prime = 5'b00101;
		10'b1001111000:	sigmoid_prime = 5'b00101;
		10'b1001111001:	sigmoid_prime = 5'b00110;
		10'b1001111010:	sigmoid_prime = 5'b00110;
		10'b1001111011:	sigmoid_prime = 5'b00110;
		10'b1001111100:	sigmoid_prime = 5'b00110;
		10'b1001111101:	sigmoid_prime = 5'b00110;
		10'b1001111110:	sigmoid_prime = 5'b00110;
		10'b1001111111:	sigmoid_prime = 5'b00110;
		10'b1010000000:	sigmoid_prime = 5'b00110;
		10'b1010000001:	sigmoid_prime = 5'b00110;
		10'b1010000010:	sigmoid_prime = 5'b00110;
		10'b1010000011:	sigmoid_prime = 5'b00110;
		10'b1010000100:	sigmoid_prime = 5'b00110;
		10'b1010000101:	sigmoid_prime = 5'b00110;
		10'b1010000110:	sigmoid_prime = 5'b00110;
		10'b1010000111:	sigmoid_prime = 5'b00110;
		10'b1010001000:	sigmoid_prime = 5'b00110;
		10'b1010001001:	sigmoid_prime = 5'b00110;
		10'b1010001010:	sigmoid_prime = 5'b00110;
		10'b1010001011:	sigmoid_prime = 5'b00110;
		10'b1010001100:	sigmoid_prime = 5'b00110;
		10'b1010001101:	sigmoid_prime = 5'b00110;
		10'b1010001110:	sigmoid_prime = 5'b00110;
		10'b1010001111:	sigmoid_prime = 5'b00110;
		10'b1010010000:	sigmoid_prime = 5'b00110;
		10'b1010010001:	sigmoid_prime = 5'b00111;
		10'b1010010010:	sigmoid_prime = 5'b00111;
		10'b1010010011:	sigmoid_prime = 5'b00111;
		10'b1010010100:	sigmoid_prime = 5'b00111;
		10'b1010010101:	sigmoid_prime = 5'b00111;
		10'b1010010110:	sigmoid_prime = 5'b00111;
		10'b1010010111:	sigmoid_prime = 5'b00111;
		10'b1010011000:	sigmoid_prime = 5'b00111;
		10'b1010011001:	sigmoid_prime = 5'b00111;
		10'b1010011010:	sigmoid_prime = 5'b00111;
		10'b1010011011:	sigmoid_prime = 5'b00111;
		10'b1010011100:	sigmoid_prime = 5'b00111;
		10'b1010011101:	sigmoid_prime = 5'b00111;
		10'b1010011110:	sigmoid_prime = 5'b00111;
		10'b1010011111:	sigmoid_prime = 5'b00111;
		10'b1010100000:	sigmoid_prime = 5'b00111;
		10'b1010100001:	sigmoid_prime = 5'b00111;
		10'b1010100010:	sigmoid_prime = 5'b00111;
		10'b1010100011:	sigmoid_prime = 5'b00111;
		10'b1010100100:	sigmoid_prime = 5'b00111;
		10'b1010100101:	sigmoid_prime = 5'b00111;
		10'b1010100110:	sigmoid_prime = 5'b01000;
		10'b1010100111:	sigmoid_prime = 5'b01000;
		10'b1010101000:	sigmoid_prime = 5'b01000;
		10'b1010101001:	sigmoid_prime = 5'b01000;
		10'b1010101010:	sigmoid_prime = 5'b01000;
		10'b1010101011:	sigmoid_prime = 5'b01000;
		10'b1010101100:	sigmoid_prime = 5'b01000;
		10'b1010101101:	sigmoid_prime = 5'b01000;
		10'b1010101110:	sigmoid_prime = 5'b01000;
		10'b1010101111:	sigmoid_prime = 5'b01000;
		10'b1010110000:	sigmoid_prime = 5'b01000;
		10'b1010110001:	sigmoid_prime = 5'b01000;
		10'b1010110010:	sigmoid_prime = 5'b01000;
		10'b1010110011:	sigmoid_prime = 5'b01000;
		10'b1010110100:	sigmoid_prime = 5'b01000;
		10'b1010110101:	sigmoid_prime = 5'b01000;
		10'b1010110110:	sigmoid_prime = 5'b01000;
		10'b1010110111:	sigmoid_prime = 5'b01000;
		10'b1010111000:	sigmoid_prime = 5'b01001;
		10'b1010111001:	sigmoid_prime = 5'b01001;
		10'b1010111010:	sigmoid_prime = 5'b01001;
		10'b1010111011:	sigmoid_prime = 5'b01001;
		10'b1010111100:	sigmoid_prime = 5'b01001;
		10'b1010111101:	sigmoid_prime = 5'b01001;
		10'b1010111110:	sigmoid_prime = 5'b01001;
		10'b1010111111:	sigmoid_prime = 5'b01001;
		10'b1011000000:	sigmoid_prime = 5'b01001;
		10'b1011000001:	sigmoid_prime = 5'b01001;
		10'b1011000010:	sigmoid_prime = 5'b01001;
		10'b1011000011:	sigmoid_prime = 5'b01001;
		10'b1011000100:	sigmoid_prime = 5'b01001;
		10'b1011000101:	sigmoid_prime = 5'b01001;
		10'b1011000110:	sigmoid_prime = 5'b01001;
		10'b1011000111:	sigmoid_prime = 5'b01001;
		10'b1011001000:	sigmoid_prime = 5'b01001;
		10'b1011001001:	sigmoid_prime = 5'b01010;
		10'b1011001010:	sigmoid_prime = 5'b01010;
		10'b1011001011:	sigmoid_prime = 5'b01010;
		10'b1011001100:	sigmoid_prime = 5'b01010;
		10'b1011001101:	sigmoid_prime = 5'b01010;
		10'b1011001110:	sigmoid_prime = 5'b01010;
		10'b1011001111:	sigmoid_prime = 5'b01010;
		10'b1011010000:	sigmoid_prime = 5'b01010;
		10'b1011010001:	sigmoid_prime = 5'b01010;
		10'b1011010010:	sigmoid_prime = 5'b01010;
		10'b1011010011:	sigmoid_prime = 5'b01010;
		10'b1011010100:	sigmoid_prime = 5'b01010;
		10'b1011010101:	sigmoid_prime = 5'b01010;
		10'b1011010110:	sigmoid_prime = 5'b01010;
		10'b1011010111:	sigmoid_prime = 5'b01010;
		10'b1011011000:	sigmoid_prime = 5'b01010;
		10'b1011011001:	sigmoid_prime = 5'b01011;
		10'b1011011010:	sigmoid_prime = 5'b01011;
		10'b1011011011:	sigmoid_prime = 5'b01011;
		10'b1011011100:	sigmoid_prime = 5'b01011;
		10'b1011011101:	sigmoid_prime = 5'b01011;
		10'b1011011110:	sigmoid_prime = 5'b01011;
		10'b1011011111:	sigmoid_prime = 5'b01011;
		10'b1011100000:	sigmoid_prime = 5'b01011;
		10'b1011100001:	sigmoid_prime = 5'b01011;
		10'b1011100010:	sigmoid_prime = 5'b01011;
		10'b1011100011:	sigmoid_prime = 5'b01011;
		10'b1011100100:	sigmoid_prime = 5'b01011;
		10'b1011100101:	sigmoid_prime = 5'b01011;
		10'b1011100110:	sigmoid_prime = 5'b01011;
		10'b1011100111:	sigmoid_prime = 5'b01100;
		10'b1011101000:	sigmoid_prime = 5'b01100;
		10'b1011101001:	sigmoid_prime = 5'b01100;
		10'b1011101010:	sigmoid_prime = 5'b01100;
		10'b1011101011:	sigmoid_prime = 5'b01100;
		10'b1011101100:	sigmoid_prime = 5'b01100;
		10'b1011101101:	sigmoid_prime = 5'b01100;
		10'b1011101110:	sigmoid_prime = 5'b01100;
		10'b1011101111:	sigmoid_prime = 5'b01100;
		10'b1011110000:	sigmoid_prime = 5'b01100;
		10'b1011110001:	sigmoid_prime = 5'b01100;
		10'b1011110010:	sigmoid_prime = 5'b01100;
		10'b1011110011:	sigmoid_prime = 5'b01100;
		10'b1011110100:	sigmoid_prime = 5'b01101;
		10'b1011110101:	sigmoid_prime = 5'b01101;
		10'b1011110110:	sigmoid_prime = 5'b01101;
		10'b1011110111:	sigmoid_prime = 5'b01101;
		10'b1011111000:	sigmoid_prime = 5'b01101;
		10'b1011111001:	sigmoid_prime = 5'b01101;
		10'b1011111010:	sigmoid_prime = 5'b01101;
		10'b1011111011:	sigmoid_prime = 5'b01101;
		10'b1011111100:	sigmoid_prime = 5'b01101;
		10'b1011111101:	sigmoid_prime = 5'b01101;
		10'b1011111110:	sigmoid_prime = 5'b01101;
		10'b1011111111:	sigmoid_prime = 5'b01101;
		10'b1100000000:	sigmoid_prime = 5'b01101;
		10'b1100000001:	sigmoid_prime = 5'b01110;
		10'b1100000010:	sigmoid_prime = 5'b01110;
		10'b1100000011:	sigmoid_prime = 5'b01110;
		10'b1100000100:	sigmoid_prime = 5'b01110;
		10'b1100000101:	sigmoid_prime = 5'b01110;
		10'b1100000110:	sigmoid_prime = 5'b01110;
		10'b1100000111:	sigmoid_prime = 5'b01110;
		10'b1100001000:	sigmoid_prime = 5'b01110;
		10'b1100001001:	sigmoid_prime = 5'b01110;
		10'b1100001010:	sigmoid_prime = 5'b01110;
		10'b1100001011:	sigmoid_prime = 5'b01110;
		10'b1100001100:	sigmoid_prime = 5'b01110;
		10'b1100001101:	sigmoid_prime = 5'b01111;
		10'b1100001110:	sigmoid_prime = 5'b01111;
		10'b1100001111:	sigmoid_prime = 5'b01111;
		10'b1100010000:	sigmoid_prime = 5'b01111;
		10'b1100010001:	sigmoid_prime = 5'b01111;
		10'b1100010010:	sigmoid_prime = 5'b01111;
		10'b1100010011:	sigmoid_prime = 5'b01111;
		10'b1100010100:	sigmoid_prime = 5'b01111;
		10'b1100010101:	sigmoid_prime = 5'b01111;
		10'b1100010110:	sigmoid_prime = 5'b01111;
		10'b1100010111:	sigmoid_prime = 5'b01111;
		10'b1100011000:	sigmoid_prime = 5'b01111;
		10'b1100011001:	sigmoid_prime = 5'b10000;
		10'b1100011010:	sigmoid_prime = 5'b10000;
		10'b1100011011:	sigmoid_prime = 5'b10000;
		10'b1100011100:	sigmoid_prime = 5'b10000;
		10'b1100011101:	sigmoid_prime = 5'b10000;
		10'b1100011110:	sigmoid_prime = 5'b10000;
		10'b1100011111:	sigmoid_prime = 5'b10000;
		10'b1100100000:	sigmoid_prime = 5'b10000;
		10'b1100100001:	sigmoid_prime = 5'b10000;
		10'b1100100010:	sigmoid_prime = 5'b10000;
		10'b1100100011:	sigmoid_prime = 5'b10000;
		10'b1100100100:	sigmoid_prime = 5'b10001;
		10'b1100100101:	sigmoid_prime = 5'b10001;
		10'b1100100110:	sigmoid_prime = 5'b10001;
		10'b1100100111:	sigmoid_prime = 5'b10001;
		10'b1100101000:	sigmoid_prime = 5'b10001;
		10'b1100101001:	sigmoid_prime = 5'b10001;
		10'b1100101010:	sigmoid_prime = 5'b10001;
		10'b1100101011:	sigmoid_prime = 5'b10001;
		10'b1100101100:	sigmoid_prime = 5'b10001;
		10'b1100101101:	sigmoid_prime = 5'b10001;
		10'b1100101110:	sigmoid_prime = 5'b10001;
		10'b1100101111:	sigmoid_prime = 5'b10010;
		10'b1100110000:	sigmoid_prime = 5'b10010;
		10'b1100110001:	sigmoid_prime = 5'b10010;
		10'b1100110010:	sigmoid_prime = 5'b10010;
		10'b1100110011:	sigmoid_prime = 5'b10010;
		10'b1100110100:	sigmoid_prime = 5'b10010;
		10'b1100110101:	sigmoid_prime = 5'b10010;
		10'b1100110110:	sigmoid_prime = 5'b10010;
		10'b1100110111:	sigmoid_prime = 5'b10010;
		10'b1100111000:	sigmoid_prime = 5'b10010;
		10'b1100111001:	sigmoid_prime = 5'b10010;
		10'b1100111010:	sigmoid_prime = 5'b10011;
		10'b1100111011:	sigmoid_prime = 5'b10011;
		10'b1100111100:	sigmoid_prime = 5'b10011;
		10'b1100111101:	sigmoid_prime = 5'b10011;
		10'b1100111110:	sigmoid_prime = 5'b10011;
		10'b1100111111:	sigmoid_prime = 5'b10011;
		10'b1101000000:	sigmoid_prime = 5'b10011;
		10'b1101000001:	sigmoid_prime = 5'b10011;
		10'b1101000010:	sigmoid_prime = 5'b10011;
		10'b1101000011:	sigmoid_prime = 5'b10011;
		10'b1101000100:	sigmoid_prime = 5'b10011;
		10'b1101000101:	sigmoid_prime = 5'b10100;
		10'b1101000110:	sigmoid_prime = 5'b10100;
		10'b1101000111:	sigmoid_prime = 5'b10100;
		10'b1101001000:	sigmoid_prime = 5'b10100;
		10'b1101001001:	sigmoid_prime = 5'b10100;
		10'b1101001010:	sigmoid_prime = 5'b10100;
		10'b1101001011:	sigmoid_prime = 5'b10100;
		10'b1101001100:	sigmoid_prime = 5'b10100;
		10'b1101001101:	sigmoid_prime = 5'b10100;
		10'b1101001110:	sigmoid_prime = 5'b10100;
		10'b1101001111:	sigmoid_prime = 5'b10101;
		10'b1101010000:	sigmoid_prime = 5'b10101;
		10'b1101010001:	sigmoid_prime = 5'b10101;
		10'b1101010010:	sigmoid_prime = 5'b10101;
		10'b1101010011:	sigmoid_prime = 5'b10101;
		10'b1101010100:	sigmoid_prime = 5'b10101;
		10'b1101010101:	sigmoid_prime = 5'b10101;
		10'b1101010110:	sigmoid_prime = 5'b10101;
		10'b1101010111:	sigmoid_prime = 5'b10101;
		10'b1101011000:	sigmoid_prime = 5'b10101;
		10'b1101011001:	sigmoid_prime = 5'b10101;
		10'b1101011010:	sigmoid_prime = 5'b10110;
		10'b1101011011:	sigmoid_prime = 5'b10110;
		10'b1101011100:	sigmoid_prime = 5'b10110;
		10'b1101011101:	sigmoid_prime = 5'b10110;
		10'b1101011110:	sigmoid_prime = 5'b10110;
		10'b1101011111:	sigmoid_prime = 5'b10110;
		10'b1101100000:	sigmoid_prime = 5'b10110;
		10'b1101100001:	sigmoid_prime = 5'b10110;
		10'b1101100010:	sigmoid_prime = 5'b10110;
		10'b1101100011:	sigmoid_prime = 5'b10110;
		10'b1101100100:	sigmoid_prime = 5'b10111;
		10'b1101100101:	sigmoid_prime = 5'b10111;
		10'b1101100110:	sigmoid_prime = 5'b10111;
		10'b1101100111:	sigmoid_prime = 5'b10111;
		10'b1101101000:	sigmoid_prime = 5'b10111;
		10'b1101101001:	sigmoid_prime = 5'b10111;
		10'b1101101010:	sigmoid_prime = 5'b10111;
		10'b1101101011:	sigmoid_prime = 5'b10111;
		10'b1101101100:	sigmoid_prime = 5'b10111;
		10'b1101101101:	sigmoid_prime = 5'b10111;
		10'b1101101110:	sigmoid_prime = 5'b10111;
		10'b1101101111:	sigmoid_prime = 5'b11000;
		10'b1101110000:	sigmoid_prime = 5'b11000;
		10'b1101110001:	sigmoid_prime = 5'b11000;
		10'b1101110010:	sigmoid_prime = 5'b11000;
		10'b1101110011:	sigmoid_prime = 5'b11000;
		10'b1101110100:	sigmoid_prime = 5'b11000;
		10'b1101110101:	sigmoid_prime = 5'b11000;
		10'b1101110110:	sigmoid_prime = 5'b11000;
		10'b1101110111:	sigmoid_prime = 5'b11000;
		10'b1101111000:	sigmoid_prime = 5'b11000;
		10'b1101111001:	sigmoid_prime = 5'b11001;
		10'b1101111010:	sigmoid_prime = 5'b11001;
		10'b1101111011:	sigmoid_prime = 5'b11001;
		10'b1101111100:	sigmoid_prime = 5'b11001;
		10'b1101111101:	sigmoid_prime = 5'b11001;
		10'b1101111110:	sigmoid_prime = 5'b11001;
		10'b1101111111:	sigmoid_prime = 5'b11001;
		10'b1110000000:	sigmoid_prime = 5'b11001;
		10'b1110000001:	sigmoid_prime = 5'b11001;
		10'b1110000010:	sigmoid_prime = 5'b11001;
		10'b1110000011:	sigmoid_prime = 5'b11001;
		10'b1110000100:	sigmoid_prime = 5'b11010;
		10'b1110000101:	sigmoid_prime = 5'b11010;
		10'b1110000110:	sigmoid_prime = 5'b11010;
		10'b1110000111:	sigmoid_prime = 5'b11010;
		10'b1110001000:	sigmoid_prime = 5'b11010;
		10'b1110001001:	sigmoid_prime = 5'b11010;
		10'b1110001010:	sigmoid_prime = 5'b11010;
		10'b1110001011:	sigmoid_prime = 5'b11010;
		10'b1110001100:	sigmoid_prime = 5'b11010;
		10'b1110001101:	sigmoid_prime = 5'b11010;
		10'b1110001110:	sigmoid_prime = 5'b11010;
		10'b1110001111:	sigmoid_prime = 5'b11010;
		10'b1110010000:	sigmoid_prime = 5'b11011;
		10'b1110010001:	sigmoid_prime = 5'b11011;
		10'b1110010010:	sigmoid_prime = 5'b11011;
		10'b1110010011:	sigmoid_prime = 5'b11011;
		10'b1110010100:	sigmoid_prime = 5'b11011;
		10'b1110010101:	sigmoid_prime = 5'b11011;
		10'b1110010110:	sigmoid_prime = 5'b11011;
		10'b1110010111:	sigmoid_prime = 5'b11011;
		10'b1110011000:	sigmoid_prime = 5'b11011;
		10'b1110011001:	sigmoid_prime = 5'b11011;
		10'b1110011010:	sigmoid_prime = 5'b11011;
		10'b1110011011:	sigmoid_prime = 5'b11011;
		10'b1110011100:	sigmoid_prime = 5'b11100;
		10'b1110011101:	sigmoid_prime = 5'b11100;
		10'b1110011110:	sigmoid_prime = 5'b11100;
		10'b1110011111:	sigmoid_prime = 5'b11100;
		10'b1110100000:	sigmoid_prime = 5'b11100;
		10'b1110100001:	sigmoid_prime = 5'b11100;
		10'b1110100010:	sigmoid_prime = 5'b11100;
		10'b1110100011:	sigmoid_prime = 5'b11100;
		10'b1110100100:	sigmoid_prime = 5'b11100;
		10'b1110100101:	sigmoid_prime = 5'b11100;
		10'b1110100110:	sigmoid_prime = 5'b11100;
		10'b1110100111:	sigmoid_prime = 5'b11100;
		10'b1110101000:	sigmoid_prime = 5'b11100;
		10'b1110101001:	sigmoid_prime = 5'b11101;
		10'b1110101010:	sigmoid_prime = 5'b11101;
		10'b1110101011:	sigmoid_prime = 5'b11101;
		10'b1110101100:	sigmoid_prime = 5'b11101;
		10'b1110101101:	sigmoid_prime = 5'b11101;
		10'b1110101110:	sigmoid_prime = 5'b11101;
		10'b1110101111:	sigmoid_prime = 5'b11101;
		10'b1110110000:	sigmoid_prime = 5'b11101;
		10'b1110110001:	sigmoid_prime = 5'b11101;
		10'b1110110010:	sigmoid_prime = 5'b11101;
		10'b1110110011:	sigmoid_prime = 5'b11101;
		10'b1110110100:	sigmoid_prime = 5'b11101;
		10'b1110110101:	sigmoid_prime = 5'b11101;
		10'b1110110110:	sigmoid_prime = 5'b11101;
		10'b1110110111:	sigmoid_prime = 5'b11110;
		10'b1110111000:	sigmoid_prime = 5'b11110;
		10'b1110111001:	sigmoid_prime = 5'b11110;
		10'b1110111010:	sigmoid_prime = 5'b11110;
		10'b1110111011:	sigmoid_prime = 5'b11110;
		10'b1110111100:	sigmoid_prime = 5'b11110;
		10'b1110111101:	sigmoid_prime = 5'b11110;
		10'b1110111110:	sigmoid_prime = 5'b11110;
		10'b1110111111:	sigmoid_prime = 5'b11110;
		10'b1111000000:	sigmoid_prime = 5'b11110;
		10'b1111000001:	sigmoid_prime = 5'b11110;
		10'b1111000010:	sigmoid_prime = 5'b11110;
		10'b1111000011:	sigmoid_prime = 5'b11110;
		10'b1111000100:	sigmoid_prime = 5'b11110;
		10'b1111000101:	sigmoid_prime = 5'b11110;
		10'b1111000110:	sigmoid_prime = 5'b11110;
		10'b1111000111:	sigmoid_prime = 5'b11110;
		10'b1111001000:	sigmoid_prime = 5'b11111;
		10'b1111001001:	sigmoid_prime = 5'b11111;
		10'b1111001010:	sigmoid_prime = 5'b11111;
		10'b1111001011:	sigmoid_prime = 5'b11111;
		10'b1111001100:	sigmoid_prime = 5'b11111;
		10'b1111001101:	sigmoid_prime = 5'b11111;
		10'b1111001110:	sigmoid_prime = 5'b11111;
		10'b1111001111:	sigmoid_prime = 5'b11111;
		10'b1111010000:	sigmoid_prime = 5'b11111;
		10'b1111010001:	sigmoid_prime = 5'b11111;
		10'b1111010010:	sigmoid_prime = 5'b11111;
		10'b1111010011:	sigmoid_prime = 5'b11111;
		10'b1111010100:	sigmoid_prime = 5'b11111;
		10'b1111010101:	sigmoid_prime = 5'b11111;
		10'b1111010110:	sigmoid_prime = 5'b11111;
		10'b1111010111:	sigmoid_prime = 5'b11111;
		10'b1111011000:	sigmoid_prime = 5'b11111;
		10'b1111011001:	sigmoid_prime = 5'b11111;
		10'b1111011010:	sigmoid_prime = 5'b11111;
		10'b1111011011:	sigmoid_prime = 5'b11111;
		10'b1111011100:	sigmoid_prime = 5'b11111;
		10'b1111011101:	sigmoid_prime = 5'b11111;
		10'b1111011110:	sigmoid_prime = 5'b11111;
		10'b1111011111:	sigmoid_prime = 5'b11111;
		10'b1111100000:	sigmoid_prime = 5'b11111;
		10'b1111100001:	sigmoid_prime = 5'b11111;
		10'b1111100010:	sigmoid_prime = 5'b11111;
		10'b1111100011:	sigmoid_prime = 5'b11111;
		10'b1111100100:	sigmoid_prime = 5'b11111;
		10'b1111100101:	sigmoid_prime = 5'b11111;
		10'b1111100110:	sigmoid_prime = 5'b11111;
		10'b1111100111:	sigmoid_prime = 5'b11111;
		10'b1111101000:	sigmoid_prime = 5'b11111;
		10'b1111101001:	sigmoid_prime = 5'b11111;
		10'b1111101010:	sigmoid_prime = 5'b11111;
		10'b1111101011:	sigmoid_prime = 5'b11111;
		10'b1111101100:	sigmoid_prime = 5'b11111;
		10'b1111101101:	sigmoid_prime = 5'b11111;
		10'b1111101110:	sigmoid_prime = 5'b11111;
		10'b1111101111:	sigmoid_prime = 5'b11111;
		10'b1111110000:	sigmoid_prime = 5'b11111;
		10'b1111110001:	sigmoid_prime = 5'b11111;
		10'b1111110010:	sigmoid_prime = 5'b11111;
		10'b1111110011:	sigmoid_prime = 5'b11111;
		10'b1111110100:	sigmoid_prime = 5'b11111;
		10'b1111110101:	sigmoid_prime = 5'b11111;
		10'b1111110110:	sigmoid_prime = 5'b11111;
		10'b1111110111:	sigmoid_prime = 5'b11111;
		10'b1111111000:	sigmoid_prime = 5'b11111;
		10'b1111111001:	sigmoid_prime = 5'b11111;
		10'b1111111010:	sigmoid_prime = 5'b11111;
		10'b1111111011:	sigmoid_prime = 5'b11111;
		10'b1111111100:	sigmoid_prime = 5'b11111;
		10'b1111111101:	sigmoid_prime = 5'b11111;
		10'b1111111110:	sigmoid_prime = 5'b11111;
		10'b1111111111:	sigmoid_prime = 5'b11111;
		10'b0000000000:	sigmoid_prime = 5'b11111;
		10'b0000000001:	sigmoid_prime = 5'b11111;
		10'b0000000010:	sigmoid_prime = 5'b11111;
		10'b0000000011:	sigmoid_prime = 5'b11111;
		10'b0000000100:	sigmoid_prime = 5'b11111;
		10'b0000000101:	sigmoid_prime = 5'b11111;
		10'b0000000110:	sigmoid_prime = 5'b11111;
		10'b0000000111:	sigmoid_prime = 5'b11111;
		10'b0000001000:	sigmoid_prime = 5'b11111;
		10'b0000001001:	sigmoid_prime = 5'b11111;
		10'b0000001010:	sigmoid_prime = 5'b11111;
		10'b0000001011:	sigmoid_prime = 5'b11111;
		10'b0000001100:	sigmoid_prime = 5'b11111;
		10'b0000001101:	sigmoid_prime = 5'b11111;
		10'b0000001110:	sigmoid_prime = 5'b11111;
		10'b0000001111:	sigmoid_prime = 5'b11111;
		10'b0000010000:	sigmoid_prime = 5'b11111;
		10'b0000010001:	sigmoid_prime = 5'b11111;
		10'b0000010010:	sigmoid_prime = 5'b11111;
		10'b0000010011:	sigmoid_prime = 5'b11111;
		10'b0000010100:	sigmoid_prime = 5'b11111;
		10'b0000010101:	sigmoid_prime = 5'b11111;
		10'b0000010110:	sigmoid_prime = 5'b11111;
		10'b0000010111:	sigmoid_prime = 5'b11111;
		10'b0000011000:	sigmoid_prime = 5'b11111;
		10'b0000011001:	sigmoid_prime = 5'b11111;
		10'b0000011010:	sigmoid_prime = 5'b11111;
		10'b0000011011:	sigmoid_prime = 5'b11111;
		10'b0000011100:	sigmoid_prime = 5'b11111;
		10'b0000011101:	sigmoid_prime = 5'b11111;
		10'b0000011110:	sigmoid_prime = 5'b11111;
		10'b0000011111:	sigmoid_prime = 5'b11111;
		10'b0000100000:	sigmoid_prime = 5'b11111;
		10'b0000100001:	sigmoid_prime = 5'b11111;
		10'b0000100010:	sigmoid_prime = 5'b11111;
		10'b0000100011:	sigmoid_prime = 5'b11111;
		10'b0000100100:	sigmoid_prime = 5'b11111;
		10'b0000100101:	sigmoid_prime = 5'b11111;
		10'b0000100110:	sigmoid_prime = 5'b11111;
		10'b0000100111:	sigmoid_prime = 5'b11111;
		10'b0000101000:	sigmoid_prime = 5'b11111;
		10'b0000101001:	sigmoid_prime = 5'b11111;
		10'b0000101010:	sigmoid_prime = 5'b11111;
		10'b0000101011:	sigmoid_prime = 5'b11111;
		10'b0000101100:	sigmoid_prime = 5'b11111;
		10'b0000101101:	sigmoid_prime = 5'b11111;
		10'b0000101110:	sigmoid_prime = 5'b11111;
		10'b0000101111:	sigmoid_prime = 5'b11111;
		10'b0000110000:	sigmoid_prime = 5'b11111;
		10'b0000110001:	sigmoid_prime = 5'b11111;
		10'b0000110010:	sigmoid_prime = 5'b11111;
		10'b0000110011:	sigmoid_prime = 5'b11111;
		10'b0000110100:	sigmoid_prime = 5'b11111;
		10'b0000110101:	sigmoid_prime = 5'b11111;
		10'b0000110110:	sigmoid_prime = 5'b11111;
		10'b0000110111:	sigmoid_prime = 5'b11111;
		10'b0000111000:	sigmoid_prime = 5'b11111;
		10'b0000111001:	sigmoid_prime = 5'b11110;
		10'b0000111010:	sigmoid_prime = 5'b11110;
		10'b0000111011:	sigmoid_prime = 5'b11110;
		10'b0000111100:	sigmoid_prime = 5'b11110;
		10'b0000111101:	sigmoid_prime = 5'b11110;
		10'b0000111110:	sigmoid_prime = 5'b11110;
		10'b0000111111:	sigmoid_prime = 5'b11110;
		10'b0001000000:	sigmoid_prime = 5'b11110;
		10'b0001000001:	sigmoid_prime = 5'b11110;
		10'b0001000010:	sigmoid_prime = 5'b11110;
		10'b0001000011:	sigmoid_prime = 5'b11110;
		10'b0001000100:	sigmoid_prime = 5'b11110;
		10'b0001000101:	sigmoid_prime = 5'b11110;
		10'b0001000110:	sigmoid_prime = 5'b11110;
		10'b0001000111:	sigmoid_prime = 5'b11110;
		10'b0001001000:	sigmoid_prime = 5'b11110;
		10'b0001001001:	sigmoid_prime = 5'b11110;
		10'b0001001010:	sigmoid_prime = 5'b11101;
		10'b0001001011:	sigmoid_prime = 5'b11101;
		10'b0001001100:	sigmoid_prime = 5'b11101;
		10'b0001001101:	sigmoid_prime = 5'b11101;
		10'b0001001110:	sigmoid_prime = 5'b11101;
		10'b0001001111:	sigmoid_prime = 5'b11101;
		10'b0001010000:	sigmoid_prime = 5'b11101;
		10'b0001010001:	sigmoid_prime = 5'b11101;
		10'b0001010010:	sigmoid_prime = 5'b11101;
		10'b0001010011:	sigmoid_prime = 5'b11101;
		10'b0001010100:	sigmoid_prime = 5'b11101;
		10'b0001010101:	sigmoid_prime = 5'b11101;
		10'b0001010110:	sigmoid_prime = 5'b11101;
		10'b0001010111:	sigmoid_prime = 5'b11101;
		10'b0001011000:	sigmoid_prime = 5'b11100;
		10'b0001011001:	sigmoid_prime = 5'b11100;
		10'b0001011010:	sigmoid_prime = 5'b11100;
		10'b0001011011:	sigmoid_prime = 5'b11100;
		10'b0001011100:	sigmoid_prime = 5'b11100;
		10'b0001011101:	sigmoid_prime = 5'b11100;
		10'b0001011110:	sigmoid_prime = 5'b11100;
		10'b0001011111:	sigmoid_prime = 5'b11100;
		10'b0001100000:	sigmoid_prime = 5'b11100;
		10'b0001100001:	sigmoid_prime = 5'b11100;
		10'b0001100010:	sigmoid_prime = 5'b11100;
		10'b0001100011:	sigmoid_prime = 5'b11100;
		10'b0001100100:	sigmoid_prime = 5'b11100;
		10'b0001100101:	sigmoid_prime = 5'b11011;
		10'b0001100110:	sigmoid_prime = 5'b11011;
		10'b0001100111:	sigmoid_prime = 5'b11011;
		10'b0001101000:	sigmoid_prime = 5'b11011;
		10'b0001101001:	sigmoid_prime = 5'b11011;
		10'b0001101010:	sigmoid_prime = 5'b11011;
		10'b0001101011:	sigmoid_prime = 5'b11011;
		10'b0001101100:	sigmoid_prime = 5'b11011;
		10'b0001101101:	sigmoid_prime = 5'b11011;
		10'b0001101110:	sigmoid_prime = 5'b11011;
		10'b0001101111:	sigmoid_prime = 5'b11011;
		10'b0001110000:	sigmoid_prime = 5'b11011;
		10'b0001110001:	sigmoid_prime = 5'b11010;
		10'b0001110010:	sigmoid_prime = 5'b11010;
		10'b0001110011:	sigmoid_prime = 5'b11010;
		10'b0001110100:	sigmoid_prime = 5'b11010;
		10'b0001110101:	sigmoid_prime = 5'b11010;
		10'b0001110110:	sigmoid_prime = 5'b11010;
		10'b0001110111:	sigmoid_prime = 5'b11010;
		10'b0001111000:	sigmoid_prime = 5'b11010;
		10'b0001111001:	sigmoid_prime = 5'b11010;
		10'b0001111010:	sigmoid_prime = 5'b11010;
		10'b0001111011:	sigmoid_prime = 5'b11010;
		10'b0001111100:	sigmoid_prime = 5'b11010;
		10'b0001111101:	sigmoid_prime = 5'b11001;
		10'b0001111110:	sigmoid_prime = 5'b11001;
		10'b0001111111:	sigmoid_prime = 5'b11001;
		10'b0010000000:	sigmoid_prime = 5'b11001;
		10'b0010000001:	sigmoid_prime = 5'b11001;
		10'b0010000010:	sigmoid_prime = 5'b11001;
		10'b0010000011:	sigmoid_prime = 5'b11001;
		10'b0010000100:	sigmoid_prime = 5'b11001;
		10'b0010000101:	sigmoid_prime = 5'b11001;
		10'b0010000110:	sigmoid_prime = 5'b11001;
		10'b0010000111:	sigmoid_prime = 5'b11001;
		10'b0010001000:	sigmoid_prime = 5'b11000;
		10'b0010001001:	sigmoid_prime = 5'b11000;
		10'b0010001010:	sigmoid_prime = 5'b11000;
		10'b0010001011:	sigmoid_prime = 5'b11000;
		10'b0010001100:	sigmoid_prime = 5'b11000;
		10'b0010001101:	sigmoid_prime = 5'b11000;
		10'b0010001110:	sigmoid_prime = 5'b11000;
		10'b0010001111:	sigmoid_prime = 5'b11000;
		10'b0010010000:	sigmoid_prime = 5'b11000;
		10'b0010010001:	sigmoid_prime = 5'b11000;
		10'b0010010010:	sigmoid_prime = 5'b10111;
		10'b0010010011:	sigmoid_prime = 5'b10111;
		10'b0010010100:	sigmoid_prime = 5'b10111;
		10'b0010010101:	sigmoid_prime = 5'b10111;
		10'b0010010110:	sigmoid_prime = 5'b10111;
		10'b0010010111:	sigmoid_prime = 5'b10111;
		10'b0010011000:	sigmoid_prime = 5'b10111;
		10'b0010011001:	sigmoid_prime = 5'b10111;
		10'b0010011010:	sigmoid_prime = 5'b10111;
		10'b0010011011:	sigmoid_prime = 5'b10111;
		10'b0010011100:	sigmoid_prime = 5'b10111;
		10'b0010011101:	sigmoid_prime = 5'b10110;
		10'b0010011110:	sigmoid_prime = 5'b10110;
		10'b0010011111:	sigmoid_prime = 5'b10110;
		10'b0010100000:	sigmoid_prime = 5'b10110;
		10'b0010100001:	sigmoid_prime = 5'b10110;
		10'b0010100010:	sigmoid_prime = 5'b10110;
		10'b0010100011:	sigmoid_prime = 5'b10110;
		10'b0010100100:	sigmoid_prime = 5'b10110;
		10'b0010100101:	sigmoid_prime = 5'b10110;
		10'b0010100110:	sigmoid_prime = 5'b10110;
		10'b0010100111:	sigmoid_prime = 5'b10101;
		10'b0010101000:	sigmoid_prime = 5'b10101;
		10'b0010101001:	sigmoid_prime = 5'b10101;
		10'b0010101010:	sigmoid_prime = 5'b10101;
		10'b0010101011:	sigmoid_prime = 5'b10101;
		10'b0010101100:	sigmoid_prime = 5'b10101;
		10'b0010101101:	sigmoid_prime = 5'b10101;
		10'b0010101110:	sigmoid_prime = 5'b10101;
		10'b0010101111:	sigmoid_prime = 5'b10101;
		10'b0010110000:	sigmoid_prime = 5'b10101;
		10'b0010110001:	sigmoid_prime = 5'b10101;
		10'b0010110010:	sigmoid_prime = 5'b10100;
		10'b0010110011:	sigmoid_prime = 5'b10100;
		10'b0010110100:	sigmoid_prime = 5'b10100;
		10'b0010110101:	sigmoid_prime = 5'b10100;
		10'b0010110110:	sigmoid_prime = 5'b10100;
		10'b0010110111:	sigmoid_prime = 5'b10100;
		10'b0010111000:	sigmoid_prime = 5'b10100;
		10'b0010111001:	sigmoid_prime = 5'b10100;
		10'b0010111010:	sigmoid_prime = 5'b10100;
		10'b0010111011:	sigmoid_prime = 5'b10100;
		10'b0010111100:	sigmoid_prime = 5'b10011;
		10'b0010111101:	sigmoid_prime = 5'b10011;
		10'b0010111110:	sigmoid_prime = 5'b10011;
		10'b0010111111:	sigmoid_prime = 5'b10011;
		10'b0011000000:	sigmoid_prime = 5'b10011;
		10'b0011000001:	sigmoid_prime = 5'b10011;
		10'b0011000010:	sigmoid_prime = 5'b10011;
		10'b0011000011:	sigmoid_prime = 5'b10011;
		10'b0011000100:	sigmoid_prime = 5'b10011;
		10'b0011000101:	sigmoid_prime = 5'b10011;
		10'b0011000110:	sigmoid_prime = 5'b10011;
		10'b0011000111:	sigmoid_prime = 5'b10010;
		10'b0011001000:	sigmoid_prime = 5'b10010;
		10'b0011001001:	sigmoid_prime = 5'b10010;
		10'b0011001010:	sigmoid_prime = 5'b10010;
		10'b0011001011:	sigmoid_prime = 5'b10010;
		10'b0011001100:	sigmoid_prime = 5'b10010;
		10'b0011001101:	sigmoid_prime = 5'b10010;
		10'b0011001110:	sigmoid_prime = 5'b10010;
		10'b0011001111:	sigmoid_prime = 5'b10010;
		10'b0011010000:	sigmoid_prime = 5'b10010;
		10'b0011010001:	sigmoid_prime = 5'b10010;
		10'b0011010010:	sigmoid_prime = 5'b10001;
		10'b0011010011:	sigmoid_prime = 5'b10001;
		10'b0011010100:	sigmoid_prime = 5'b10001;
		10'b0011010101:	sigmoid_prime = 5'b10001;
		10'b0011010110:	sigmoid_prime = 5'b10001;
		10'b0011010111:	sigmoid_prime = 5'b10001;
		10'b0011011000:	sigmoid_prime = 5'b10001;
		10'b0011011001:	sigmoid_prime = 5'b10001;
		10'b0011011010:	sigmoid_prime = 5'b10001;
		10'b0011011011:	sigmoid_prime = 5'b10001;
		10'b0011011100:	sigmoid_prime = 5'b10001;
		10'b0011011101:	sigmoid_prime = 5'b10000;
		10'b0011011110:	sigmoid_prime = 5'b10000;
		10'b0011011111:	sigmoid_prime = 5'b10000;
		10'b0011100000:	sigmoid_prime = 5'b10000;
		10'b0011100001:	sigmoid_prime = 5'b10000;
		10'b0011100010:	sigmoid_prime = 5'b10000;
		10'b0011100011:	sigmoid_prime = 5'b10000;
		10'b0011100100:	sigmoid_prime = 5'b10000;
		10'b0011100101:	sigmoid_prime = 5'b10000;
		10'b0011100110:	sigmoid_prime = 5'b10000;
		10'b0011100111:	sigmoid_prime = 5'b10000;
		10'b0011101000:	sigmoid_prime = 5'b01111;
		10'b0011101001:	sigmoid_prime = 5'b01111;
		10'b0011101010:	sigmoid_prime = 5'b01111;
		10'b0011101011:	sigmoid_prime = 5'b01111;
		10'b0011101100:	sigmoid_prime = 5'b01111;
		10'b0011101101:	sigmoid_prime = 5'b01111;
		10'b0011101110:	sigmoid_prime = 5'b01111;
		10'b0011101111:	sigmoid_prime = 5'b01111;
		10'b0011110000:	sigmoid_prime = 5'b01111;
		10'b0011110001:	sigmoid_prime = 5'b01111;
		10'b0011110010:	sigmoid_prime = 5'b01111;
		10'b0011110011:	sigmoid_prime = 5'b01111;
		10'b0011110100:	sigmoid_prime = 5'b01110;
		10'b0011110101:	sigmoid_prime = 5'b01110;
		10'b0011110110:	sigmoid_prime = 5'b01110;
		10'b0011110111:	sigmoid_prime = 5'b01110;
		10'b0011111000:	sigmoid_prime = 5'b01110;
		10'b0011111001:	sigmoid_prime = 5'b01110;
		10'b0011111010:	sigmoid_prime = 5'b01110;
		10'b0011111011:	sigmoid_prime = 5'b01110;
		10'b0011111100:	sigmoid_prime = 5'b01110;
		10'b0011111101:	sigmoid_prime = 5'b01110;
		10'b0011111110:	sigmoid_prime = 5'b01110;
		10'b0011111111:	sigmoid_prime = 5'b01110;
		10'b0100000000:	sigmoid_prime = 5'b01101;
		10'b0100000001:	sigmoid_prime = 5'b01101;
		10'b0100000010:	sigmoid_prime = 5'b01101;
		10'b0100000011:	sigmoid_prime = 5'b01101;
		10'b0100000100:	sigmoid_prime = 5'b01101;
		10'b0100000101:	sigmoid_prime = 5'b01101;
		10'b0100000110:	sigmoid_prime = 5'b01101;
		10'b0100000111:	sigmoid_prime = 5'b01101;
		10'b0100001000:	sigmoid_prime = 5'b01101;
		10'b0100001001:	sigmoid_prime = 5'b01101;
		10'b0100001010:	sigmoid_prime = 5'b01101;
		10'b0100001011:	sigmoid_prime = 5'b01101;
		10'b0100001100:	sigmoid_prime = 5'b01101;
		10'b0100001101:	sigmoid_prime = 5'b01100;
		10'b0100001110:	sigmoid_prime = 5'b01100;
		10'b0100001111:	sigmoid_prime = 5'b01100;
		10'b0100010000:	sigmoid_prime = 5'b01100;
		10'b0100010001:	sigmoid_prime = 5'b01100;
		10'b0100010010:	sigmoid_prime = 5'b01100;
		10'b0100010011:	sigmoid_prime = 5'b01100;
		10'b0100010100:	sigmoid_prime = 5'b01100;
		10'b0100010101:	sigmoid_prime = 5'b01100;
		10'b0100010110:	sigmoid_prime = 5'b01100;
		10'b0100010111:	sigmoid_prime = 5'b01100;
		10'b0100011000:	sigmoid_prime = 5'b01100;
		10'b0100011001:	sigmoid_prime = 5'b01100;
		10'b0100011010:	sigmoid_prime = 5'b01011;
		10'b0100011011:	sigmoid_prime = 5'b01011;
		10'b0100011100:	sigmoid_prime = 5'b01011;
		10'b0100011101:	sigmoid_prime = 5'b01011;
		10'b0100011110:	sigmoid_prime = 5'b01011;
		10'b0100011111:	sigmoid_prime = 5'b01011;
		10'b0100100000:	sigmoid_prime = 5'b01011;
		10'b0100100001:	sigmoid_prime = 5'b01011;
		10'b0100100010:	sigmoid_prime = 5'b01011;
		10'b0100100011:	sigmoid_prime = 5'b01011;
		10'b0100100100:	sigmoid_prime = 5'b01011;
		10'b0100100101:	sigmoid_prime = 5'b01011;
		10'b0100100110:	sigmoid_prime = 5'b01011;
		10'b0100100111:	sigmoid_prime = 5'b01011;
		10'b0100101000:	sigmoid_prime = 5'b01010;
		10'b0100101001:	sigmoid_prime = 5'b01010;
		10'b0100101010:	sigmoid_prime = 5'b01010;
		10'b0100101011:	sigmoid_prime = 5'b01010;
		10'b0100101100:	sigmoid_prime = 5'b01010;
		10'b0100101101:	sigmoid_prime = 5'b01010;
		10'b0100101110:	sigmoid_prime = 5'b01010;
		10'b0100101111:	sigmoid_prime = 5'b01010;
		10'b0100110000:	sigmoid_prime = 5'b01010;
		10'b0100110001:	sigmoid_prime = 5'b01010;
		10'b0100110010:	sigmoid_prime = 5'b01010;
		10'b0100110011:	sigmoid_prime = 5'b01010;
		10'b0100110100:	sigmoid_prime = 5'b01010;
		10'b0100110101:	sigmoid_prime = 5'b01010;
		10'b0100110110:	sigmoid_prime = 5'b01010;
		10'b0100110111:	sigmoid_prime = 5'b01010;
		10'b0100111000:	sigmoid_prime = 5'b01001;
		10'b0100111001:	sigmoid_prime = 5'b01001;
		10'b0100111010:	sigmoid_prime = 5'b01001;
		10'b0100111011:	sigmoid_prime = 5'b01001;
		10'b0100111100:	sigmoid_prime = 5'b01001;
		10'b0100111101:	sigmoid_prime = 5'b01001;
		10'b0100111110:	sigmoid_prime = 5'b01001;
		10'b0100111111:	sigmoid_prime = 5'b01001;
		10'b0101000000:	sigmoid_prime = 5'b01001;
		10'b0101000001:	sigmoid_prime = 5'b01001;
		10'b0101000010:	sigmoid_prime = 5'b01001;
		10'b0101000011:	sigmoid_prime = 5'b01001;
		10'b0101000100:	sigmoid_prime = 5'b01001;
		10'b0101000101:	sigmoid_prime = 5'b01001;
		10'b0101000110:	sigmoid_prime = 5'b01001;
		10'b0101000111:	sigmoid_prime = 5'b01001;
		10'b0101001000:	sigmoid_prime = 5'b01001;
		10'b0101001001:	sigmoid_prime = 5'b01000;
		10'b0101001010:	sigmoid_prime = 5'b01000;
		10'b0101001011:	sigmoid_prime = 5'b01000;
		10'b0101001100:	sigmoid_prime = 5'b01000;
		10'b0101001101:	sigmoid_prime = 5'b01000;
		10'b0101001110:	sigmoid_prime = 5'b01000;
		10'b0101001111:	sigmoid_prime = 5'b01000;
		10'b0101010000:	sigmoid_prime = 5'b01000;
		10'b0101010001:	sigmoid_prime = 5'b01000;
		10'b0101010010:	sigmoid_prime = 5'b01000;
		10'b0101010011:	sigmoid_prime = 5'b01000;
		10'b0101010100:	sigmoid_prime = 5'b01000;
		10'b0101010101:	sigmoid_prime = 5'b01000;
		10'b0101010110:	sigmoid_prime = 5'b01000;
		10'b0101010111:	sigmoid_prime = 5'b01000;
		10'b0101011000:	sigmoid_prime = 5'b01000;
		10'b0101011001:	sigmoid_prime = 5'b01000;
		10'b0101011010:	sigmoid_prime = 5'b01000;
		10'b0101011011:	sigmoid_prime = 5'b00111;
		10'b0101011100:	sigmoid_prime = 5'b00111;
		10'b0101011101:	sigmoid_prime = 5'b00111;
		10'b0101011110:	sigmoid_prime = 5'b00111;
		10'b0101011111:	sigmoid_prime = 5'b00111;
		10'b0101100000:	sigmoid_prime = 5'b00111;
		10'b0101100001:	sigmoid_prime = 5'b00111;
		10'b0101100010:	sigmoid_prime = 5'b00111;
		10'b0101100011:	sigmoid_prime = 5'b00111;
		10'b0101100100:	sigmoid_prime = 5'b00111;
		10'b0101100101:	sigmoid_prime = 5'b00111;
		10'b0101100110:	sigmoid_prime = 5'b00111;
		10'b0101100111:	sigmoid_prime = 5'b00111;
		10'b0101101000:	sigmoid_prime = 5'b00111;
		10'b0101101001:	sigmoid_prime = 5'b00111;
		10'b0101101010:	sigmoid_prime = 5'b00111;
		10'b0101101011:	sigmoid_prime = 5'b00111;
		10'b0101101100:	sigmoid_prime = 5'b00111;
		10'b0101101101:	sigmoid_prime = 5'b00111;
		10'b0101101110:	sigmoid_prime = 5'b00111;
		10'b0101101111:	sigmoid_prime = 5'b00111;
		10'b0101110000:	sigmoid_prime = 5'b00110;
		10'b0101110001:	sigmoid_prime = 5'b00110;
		10'b0101110010:	sigmoid_prime = 5'b00110;
		10'b0101110011:	sigmoid_prime = 5'b00110;
		10'b0101110100:	sigmoid_prime = 5'b00110;
		10'b0101110101:	sigmoid_prime = 5'b00110;
		10'b0101110110:	sigmoid_prime = 5'b00110;
		10'b0101110111:	sigmoid_prime = 5'b00110;
		10'b0101111000:	sigmoid_prime = 5'b00110;
		10'b0101111001:	sigmoid_prime = 5'b00110;
		10'b0101111010:	sigmoid_prime = 5'b00110;
		10'b0101111011:	sigmoid_prime = 5'b00110;
		10'b0101111100:	sigmoid_prime = 5'b00110;
		10'b0101111101:	sigmoid_prime = 5'b00110;
		10'b0101111110:	sigmoid_prime = 5'b00110;
		10'b0101111111:	sigmoid_prime = 5'b00110;
		10'b0110000000:	sigmoid_prime = 5'b00110;
		10'b0110000001:	sigmoid_prime = 5'b00110;
		10'b0110000010:	sigmoid_prime = 5'b00110;
		10'b0110000011:	sigmoid_prime = 5'b00110;
		10'b0110000100:	sigmoid_prime = 5'b00110;
		10'b0110000101:	sigmoid_prime = 5'b00110;
		10'b0110000110:	sigmoid_prime = 5'b00110;
		10'b0110000111:	sigmoid_prime = 5'b00110;
		10'b0110001000:	sigmoid_prime = 5'b00101;
		10'b0110001001:	sigmoid_prime = 5'b00101;
		10'b0110001010:	sigmoid_prime = 5'b00101;
		10'b0110001011:	sigmoid_prime = 5'b00101;
		10'b0110001100:	sigmoid_prime = 5'b00101;
		10'b0110001101:	sigmoid_prime = 5'b00101;
		10'b0110001110:	sigmoid_prime = 5'b00101;
		10'b0110001111:	sigmoid_prime = 5'b00101;
		10'b0110010000:	sigmoid_prime = 5'b00101;
		10'b0110010001:	sigmoid_prime = 5'b00101;
		10'b0110010010:	sigmoid_prime = 5'b00101;
		10'b0110010011:	sigmoid_prime = 5'b00101;
		10'b0110010100:	sigmoid_prime = 5'b00101;
		10'b0110010101:	sigmoid_prime = 5'b00101;
		10'b0110010110:	sigmoid_prime = 5'b00101;
		10'b0110010111:	sigmoid_prime = 5'b00101;
		10'b0110011000:	sigmoid_prime = 5'b00101;
		10'b0110011001:	sigmoid_prime = 5'b00101;
		10'b0110011010:	sigmoid_prime = 5'b00101;
		10'b0110011011:	sigmoid_prime = 5'b00101;
		10'b0110011100:	sigmoid_prime = 5'b00101;
		10'b0110011101:	sigmoid_prime = 5'b00101;
		10'b0110011110:	sigmoid_prime = 5'b00101;
		10'b0110011111:	sigmoid_prime = 5'b00101;
		10'b0110100000:	sigmoid_prime = 5'b00101;
		10'b0110100001:	sigmoid_prime = 5'b00101;
		10'b0110100010:	sigmoid_prime = 5'b00101;
		10'b0110100011:	sigmoid_prime = 5'b00101;
		10'b0110100100:	sigmoid_prime = 5'b00100;
		10'b0110100101:	sigmoid_prime = 5'b00100;
		10'b0110100110:	sigmoid_prime = 5'b00100;
		10'b0110100111:	sigmoid_prime = 5'b00100;
		10'b0110101000:	sigmoid_prime = 5'b00100;
		10'b0110101001:	sigmoid_prime = 5'b00100;
		10'b0110101010:	sigmoid_prime = 5'b00100;
		10'b0110101011:	sigmoid_prime = 5'b00100;
		10'b0110101100:	sigmoid_prime = 5'b00100;
		10'b0110101101:	sigmoid_prime = 5'b00100;
		10'b0110101110:	sigmoid_prime = 5'b00100;
		10'b0110101111:	sigmoid_prime = 5'b00100;
		10'b0110110000:	sigmoid_prime = 5'b00100;
		10'b0110110001:	sigmoid_prime = 5'b00100;
		10'b0110110010:	sigmoid_prime = 5'b00100;
		10'b0110110011:	sigmoid_prime = 5'b00100;
		10'b0110110100:	sigmoid_prime = 5'b00100;
		10'b0110110101:	sigmoid_prime = 5'b00100;
		10'b0110110110:	sigmoid_prime = 5'b00100;
		10'b0110110111:	sigmoid_prime = 5'b00100;
		10'b0110111000:	sigmoid_prime = 5'b00100;
		10'b0110111001:	sigmoid_prime = 5'b00100;
		10'b0110111010:	sigmoid_prime = 5'b00100;
		10'b0110111011:	sigmoid_prime = 5'b00100;
		10'b0110111100:	sigmoid_prime = 5'b00100;
		10'b0110111101:	sigmoid_prime = 5'b00100;
		10'b0110111110:	sigmoid_prime = 5'b00100;
		10'b0110111111:	sigmoid_prime = 5'b00100;
		10'b0111000000:	sigmoid_prime = 5'b00100;
		10'b0111000001:	sigmoid_prime = 5'b00100;
		10'b0111000010:	sigmoid_prime = 5'b00100;
		10'b0111000011:	sigmoid_prime = 5'b00100;
		10'b0111000100:	sigmoid_prime = 5'b00100;
		10'b0111000101:	sigmoid_prime = 5'b00100;
		10'b0111000110:	sigmoid_prime = 5'b00011;
		10'b0111000111:	sigmoid_prime = 5'b00011;
		10'b0111001000:	sigmoid_prime = 5'b00011;
		10'b0111001001:	sigmoid_prime = 5'b00011;
		10'b0111001010:	sigmoid_prime = 5'b00011;
		10'b0111001011:	sigmoid_prime = 5'b00011;
		10'b0111001100:	sigmoid_prime = 5'b00011;
		10'b0111001101:	sigmoid_prime = 5'b00011;
		10'b0111001110:	sigmoid_prime = 5'b00011;
		10'b0111001111:	sigmoid_prime = 5'b00011;
		10'b0111010000:	sigmoid_prime = 5'b00011;
		10'b0111010001:	sigmoid_prime = 5'b00011;
		10'b0111010010:	sigmoid_prime = 5'b00011;
		10'b0111010011:	sigmoid_prime = 5'b00011;
		10'b0111010100:	sigmoid_prime = 5'b00011;
		10'b0111010101:	sigmoid_prime = 5'b00011;
		10'b0111010110:	sigmoid_prime = 5'b00011;
		10'b0111010111:	sigmoid_prime = 5'b00011;
		10'b0111011000:	sigmoid_prime = 5'b00011;
		10'b0111011001:	sigmoid_prime = 5'b00011;
		10'b0111011010:	sigmoid_prime = 5'b00011;
		10'b0111011011:	sigmoid_prime = 5'b00011;
		10'b0111011100:	sigmoid_prime = 5'b00011;
		10'b0111011101:	sigmoid_prime = 5'b00011;
		10'b0111011110:	sigmoid_prime = 5'b00011;
		10'b0111011111:	sigmoid_prime = 5'b00011;
		10'b0111100000:	sigmoid_prime = 5'b00011;
		10'b0111100001:	sigmoid_prime = 5'b00011;
		10'b0111100010:	sigmoid_prime = 5'b00011;
		10'b0111100011:	sigmoid_prime = 5'b00011;
		10'b0111100100:	sigmoid_prime = 5'b00011;
		10'b0111100101:	sigmoid_prime = 5'b00011;
		10'b0111100110:	sigmoid_prime = 5'b00011;
		10'b0111100111:	sigmoid_prime = 5'b00011;
		10'b0111101000:	sigmoid_prime = 5'b00011;
		10'b0111101001:	sigmoid_prime = 5'b00011;
		10'b0111101010:	sigmoid_prime = 5'b00011;
		10'b0111101011:	sigmoid_prime = 5'b00011;
		10'b0111101100:	sigmoid_prime = 5'b00011;
		10'b0111101101:	sigmoid_prime = 5'b00011;
		10'b0111101110:	sigmoid_prime = 5'b00011;
		10'b0111101111:	sigmoid_prime = 5'b00011;
		10'b0111110000:	sigmoid_prime = 5'b00011;
		10'b0111110001:	sigmoid_prime = 5'b00011;
		10'b0111110010:	sigmoid_prime = 5'b00011;
		10'b0111110011:	sigmoid_prime = 5'b00010;
		10'b0111110100:	sigmoid_prime = 5'b00010;
		10'b0111110101:	sigmoid_prime = 5'b00010;
		10'b0111110110:	sigmoid_prime = 5'b00010;
		10'b0111110111:	sigmoid_prime = 5'b00010;
		10'b0111111000:	sigmoid_prime = 5'b00010;
		10'b0111111001:	sigmoid_prime = 5'b00010;
		10'b0111111010:	sigmoid_prime = 5'b00010;
		10'b0111111011:	sigmoid_prime = 5'b00010;
		10'b0111111100:	sigmoid_prime = 5'b00010;
		10'b0111111101:	sigmoid_prime = 5'b00010;
		10'b0111111110:	sigmoid_prime = 5'b00010;
		10'b0111111111:	sigmoid_prime = 5'b00010;

	endcase
endmodule
