// Activation functions using clock, i.e. act and actprime available at next posedge
// Sourya Dey, Yinan Shao, USC

// If any parameter is changed, sigmoid tables will have to be regenerated using dnn-rtl/scripts/actlut_generator.py
// To be replaced in sigmoid: parameter values, and the table portion inside the case statements. Nothing else.
// NOTHING IN RELU EVER NEEDS TO BE REPLACED, IT IS COMPLETELY PARAMETRIZED

`timescale 1ns/100ps

module relu_all #(
	parameter width = 12,
	parameter int_bits = 3,
	localparam frac_bits = width-int_bits-1
)(
	input clk,
	input signed [width-1:0] val,
	output logic [width-1:0] relu_out = '0,
	output logic [width-1:0] relu_prime_out = '0
);

	// Use raw values to mimic coding style in sigmoid
	logic [width-1:0] relu = '0;
	logic [width-1:0] relu_prime = '0;
	
	always @(posedge clk) begin	
		relu_out <= relu;
		relu_prime_out <= relu_prime;
	end
	
	always_comb begin
		relu <= (val <= 0) ? 1 : (val >= 1<<frac_bits) ? {{(int_bits+1){1'b0}},{(frac_bits){1'b1}}} : val;
		relu_prime <= ((val <= 0) || (val >= 1<<frac_bits)) ? 1 : {{(int_bits+1){1'b0}},{(frac_bits){1'b1}}};
	end
endmodule


module sigmoid_all #(
	parameter width = 12,
	parameter int_bits = 3,
	localparam frac_bits = width-int_bits-1,
	parameter maxdomain = (2**int_bits>8) ? 8 : 2**int_bits, //8 is arbitrarily chosen
	//input has to be within [-maxdomain,maxdomain). If outside this range, sigmoid is either 0 or 1
	parameter lut_size_prelim = (2**width>4096) ? 4096 : 2**width, //4096 is arbitrarily chosen
	localparam lut_size = (lut_size_prelim > 2**(frac_bits+$clog2(maxdomain)+1)) ? 2**(frac_bits+$clog2(maxdomain)+1) : lut_size_prelim //actual lut_size
	// If lut_size is > 2**(frac_bits+$clog2(maxdomain)+1)), then val[frac_bits+$clog2(maxdomain) -: $clog2(lut_size)] would be an invalid part select
	// Ideally they should not, but it could happen that maxdomain and lut_size_prelim are set from outside, so they are params, not localparams
)(
	input clk,
	input signed [width-1:0] val,
	output logic [width-1:0] sigmoid_out = '0,
	output logic [width-1:0] sigmoid_prime_out = '0
);

	logic [frac_bits-1:0] sigmoid = '0; //raw sigmoid value
	logic [frac_bits-3:0] sigmoid_prime = '0; //raw sigmoid_prime value, 2 bits less since 2 MSB in frac_part are always 00

	always @(posedge clk) begin
		sigmoid_out <= (val[width-1 : frac_bits+$clog2(maxdomain)] == 0 || &val[width-1 : frac_bits+$clog2(maxdomain)]) ? // Only calculate sigmoid for the domain val = [-maxdomain,+maxdomain). So check all MSB till there. If all 0, val<maxdomain. If all 1, val>=-maxdomain
		{{(int_bits+1){1'b0}}, sigmoid} : //If val is within [-maxdomain,+maxdomain), insert all 0s for sign and integer part (since sigmoid is always between 0 and 1) and then frac_bits sigmoid part
		(val[width-1]) ? //If val is outside the range, sigmoid will be 0 or 1 depending on sign bit
		1 : //If sign bit is 1, val is negative, so sigmoid is 0
		{{(int_bits+1){1'b0}},{(frac_bits){1'b1}}}; //If sign bit is 0, val is positive. Then sigmoid is all 1s in the fractional part, i.e. 1-2^(-frac_bits), which is the highest number possible (~=1)

		sigmoid_prime_out <= (val[width-1 : frac_bits+$clog2(maxdomain)] == 0 || &val[width-1 : frac_bits+$clog2(maxdomain)]) ? 
		{{(int_bits+3){1'b0}},sigmoid_prime} : //since 2 MSB in frac_part are always 00
		1; //If val is outside [-maxdomain,+maxdomain], sigmoid prime will always be 0
	end

	always_comb begin
	case (val[frac_bits+$clog2(maxdomain) -: $clog2(lut_size)]) //this ensures that we read exactly log(lut_size) bits as address of LUT
		
				10'b1000000000: begin sigmoid <= 7'b0000010; sigmoid_prime <= 5'b00010; end
				10'b1000000001: begin sigmoid <= 7'b0000010; sigmoid_prime <= 5'b00010; end
				10'b1000000010: begin sigmoid <= 7'b0000010; sigmoid_prime <= 5'b00010; end
				10'b1000000011: begin sigmoid <= 7'b0000010; sigmoid_prime <= 5'b00010; end
				10'b1000000100: begin sigmoid <= 7'b0000010; sigmoid_prime <= 5'b00010; end
				10'b1000000101: begin sigmoid <= 7'b0000010; sigmoid_prime <= 5'b00010; end
				10'b1000000110: begin sigmoid <= 7'b0000010; sigmoid_prime <= 5'b00010; end
				10'b1000000111: begin sigmoid <= 7'b0000010; sigmoid_prime <= 5'b00010; end
				10'b1000001000: begin sigmoid <= 7'b0000010; sigmoid_prime <= 5'b00010; end
				10'b1000001001: begin sigmoid <= 7'b0000010; sigmoid_prime <= 5'b00010; end
				10'b1000001010: begin sigmoid <= 7'b0000010; sigmoid_prime <= 5'b00010; end
				10'b1000001011: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00010; end
				10'b1000001100: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00010; end
				10'b1000001101: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00010; end
				10'b1000001110: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000001111: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000010000: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000010001: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000010010: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000010011: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000010100: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000010101: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000010110: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000010111: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000011000: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000011001: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000011010: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000011011: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000011100: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000011101: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000011110: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000011111: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000100000: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000100001: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000100010: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000100011: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000100100: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000100101: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000100110: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000100111: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000101000: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000101001: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000101010: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000101011: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000101100: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000101101: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000101110: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000101111: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000110000: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000110001: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000110010: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000110011: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000110100: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000110101: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000110110: begin sigmoid <= 7'b0000011; sigmoid_prime <= 5'b00011; end
				10'b1000110111: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00011; end
				10'b1000111000: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00011; end
				10'b1000111001: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00011; end
				10'b1000111010: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00011; end
				10'b1000111011: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1000111100: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1000111101: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1000111110: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1000111111: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001000000: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001000001: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001000010: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001000011: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001000100: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001000101: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001000110: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001000111: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001001000: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001001001: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001001010: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001001011: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001001100: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001001101: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001001110: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001001111: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001010000: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001010001: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001010010: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001010011: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001010100: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001010101: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001010110: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001010111: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001011000: begin sigmoid <= 7'b0000100; sigmoid_prime <= 5'b00100; end
				10'b1001011001: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00100; end
				10'b1001011010: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00100; end
				10'b1001011011: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00100; end
				10'b1001011100: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00100; end
				10'b1001011101: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001011110: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001011111: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001100000: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001100001: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001100010: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001100011: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001100100: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001100101: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001100110: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001100111: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001101000: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001101001: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001101010: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001101011: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001101100: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001101101: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001101110: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001101111: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001110000: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001110001: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001110010: begin sigmoid <= 7'b0000101; sigmoid_prime <= 5'b00101; end
				10'b1001110011: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00101; end
				10'b1001110100: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00101; end
				10'b1001110101: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00101; end
				10'b1001110110: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00101; end
				10'b1001110111: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00101; end
				10'b1001111000: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00101; end
				10'b1001111001: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1001111010: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1001111011: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1001111100: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1001111101: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1001111110: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1001111111: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1010000000: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1010000001: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1010000010: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1010000011: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1010000100: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1010000101: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1010000110: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1010000111: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1010001000: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1010001001: begin sigmoid <= 7'b0000110; sigmoid_prime <= 5'b00110; end
				10'b1010001010: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00110; end
				10'b1010001011: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00110; end
				10'b1010001100: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00110; end
				10'b1010001101: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00110; end
				10'b1010001110: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00110; end
				10'b1010001111: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00110; end
				10'b1010010000: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00110; end
				10'b1010010001: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00111; end
				10'b1010010010: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00111; end
				10'b1010010011: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00111; end
				10'b1010010100: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00111; end
				10'b1010010101: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00111; end
				10'b1010010110: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00111; end
				10'b1010010111: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00111; end
				10'b1010011000: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00111; end
				10'b1010011001: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00111; end
				10'b1010011010: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00111; end
				10'b1010011011: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00111; end
				10'b1010011100: begin sigmoid <= 7'b0000111; sigmoid_prime <= 5'b00111; end
				10'b1010011101: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b00111; end
				10'b1010011110: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b00111; end
				10'b1010011111: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b00111; end
				10'b1010100000: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b00111; end
				10'b1010100001: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b00111; end
				10'b1010100010: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b00111; end
				10'b1010100011: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b00111; end
				10'b1010100100: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b00111; end
				10'b1010100101: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b00111; end
				10'b1010100110: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b01000; end
				10'b1010100111: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b01000; end
				10'b1010101000: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b01000; end
				10'b1010101001: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b01000; end
				10'b1010101010: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b01000; end
				10'b1010101011: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b01000; end
				10'b1010101100: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b01000; end
				10'b1010101101: begin sigmoid <= 7'b0001000; sigmoid_prime <= 5'b01000; end
				10'b1010101110: begin sigmoid <= 7'b0001001; sigmoid_prime <= 5'b01000; end
				10'b1010101111: begin sigmoid <= 7'b0001001; sigmoid_prime <= 5'b01000; end
				10'b1010110000: begin sigmoid <= 7'b0001001; sigmoid_prime <= 5'b01000; end
				10'b1010110001: begin sigmoid <= 7'b0001001; sigmoid_prime <= 5'b01000; end
				10'b1010110010: begin sigmoid <= 7'b0001001; sigmoid_prime <= 5'b01000; end
				10'b1010110011: begin sigmoid <= 7'b0001001; sigmoid_prime <= 5'b01000; end
				10'b1010110100: begin sigmoid <= 7'b0001001; sigmoid_prime <= 5'b01000; end
				10'b1010110101: begin sigmoid <= 7'b0001001; sigmoid_prime <= 5'b01000; end
				10'b1010110110: begin sigmoid <= 7'b0001001; sigmoid_prime <= 5'b01000; end
				10'b1010110111: begin sigmoid <= 7'b0001001; sigmoid_prime <= 5'b01000; end
				10'b1010111000: begin sigmoid <= 7'b0001001; sigmoid_prime <= 5'b01001; end
				10'b1010111001: begin sigmoid <= 7'b0001001; sigmoid_prime <= 5'b01001; end
				10'b1010111010: begin sigmoid <= 7'b0001001; sigmoid_prime <= 5'b01001; end
				10'b1010111011: begin sigmoid <= 7'b0001001; sigmoid_prime <= 5'b01001; end
				10'b1010111100: begin sigmoid <= 7'b0001001; sigmoid_prime <= 5'b01001; end
				10'b1010111101: begin sigmoid <= 7'b0001010; sigmoid_prime <= 5'b01001; end
				10'b1010111110: begin sigmoid <= 7'b0001010; sigmoid_prime <= 5'b01001; end
				10'b1010111111: begin sigmoid <= 7'b0001010; sigmoid_prime <= 5'b01001; end
				10'b1011000000: begin sigmoid <= 7'b0001010; sigmoid_prime <= 5'b01001; end
				10'b1011000001: begin sigmoid <= 7'b0001010; sigmoid_prime <= 5'b01001; end
				10'b1011000010: begin sigmoid <= 7'b0001010; sigmoid_prime <= 5'b01001; end
				10'b1011000011: begin sigmoid <= 7'b0001010; sigmoid_prime <= 5'b01001; end
				10'b1011000100: begin sigmoid <= 7'b0001010; sigmoid_prime <= 5'b01001; end
				10'b1011000101: begin sigmoid <= 7'b0001010; sigmoid_prime <= 5'b01001; end
				10'b1011000110: begin sigmoid <= 7'b0001010; sigmoid_prime <= 5'b01001; end
				10'b1011000111: begin sigmoid <= 7'b0001010; sigmoid_prime <= 5'b01001; end
				10'b1011001000: begin sigmoid <= 7'b0001010; sigmoid_prime <= 5'b01001; end
				10'b1011001001: begin sigmoid <= 7'b0001010; sigmoid_prime <= 5'b01010; end
				10'b1011001010: begin sigmoid <= 7'b0001010; sigmoid_prime <= 5'b01010; end
				10'b1011001011: begin sigmoid <= 7'b0001011; sigmoid_prime <= 5'b01010; end
				10'b1011001100: begin sigmoid <= 7'b0001011; sigmoid_prime <= 5'b01010; end
				10'b1011001101: begin sigmoid <= 7'b0001011; sigmoid_prime <= 5'b01010; end
				10'b1011001110: begin sigmoid <= 7'b0001011; sigmoid_prime <= 5'b01010; end
				10'b1011001111: begin sigmoid <= 7'b0001011; sigmoid_prime <= 5'b01010; end
				10'b1011010000: begin sigmoid <= 7'b0001011; sigmoid_prime <= 5'b01010; end
				10'b1011010001: begin sigmoid <= 7'b0001011; sigmoid_prime <= 5'b01010; end
				10'b1011010010: begin sigmoid <= 7'b0001011; sigmoid_prime <= 5'b01010; end
				10'b1011010011: begin sigmoid <= 7'b0001011; sigmoid_prime <= 5'b01010; end
				10'b1011010100: begin sigmoid <= 7'b0001011; sigmoid_prime <= 5'b01010; end
				10'b1011010101: begin sigmoid <= 7'b0001011; sigmoid_prime <= 5'b01010; end
				10'b1011010110: begin sigmoid <= 7'b0001011; sigmoid_prime <= 5'b01010; end
				10'b1011010111: begin sigmoid <= 7'b0001011; sigmoid_prime <= 5'b01010; end
				10'b1011011000: begin sigmoid <= 7'b0001100; sigmoid_prime <= 5'b01010; end
				10'b1011011001: begin sigmoid <= 7'b0001100; sigmoid_prime <= 5'b01011; end
				10'b1011011010: begin sigmoid <= 7'b0001100; sigmoid_prime <= 5'b01011; end
				10'b1011011011: begin sigmoid <= 7'b0001100; sigmoid_prime <= 5'b01011; end
				10'b1011011100: begin sigmoid <= 7'b0001100; sigmoid_prime <= 5'b01011; end
				10'b1011011101: begin sigmoid <= 7'b0001100; sigmoid_prime <= 5'b01011; end
				10'b1011011110: begin sigmoid <= 7'b0001100; sigmoid_prime <= 5'b01011; end
				10'b1011011111: begin sigmoid <= 7'b0001100; sigmoid_prime <= 5'b01011; end
				10'b1011100000: begin sigmoid <= 7'b0001100; sigmoid_prime <= 5'b01011; end
				10'b1011100001: begin sigmoid <= 7'b0001100; sigmoid_prime <= 5'b01011; end
				10'b1011100010: begin sigmoid <= 7'b0001100; sigmoid_prime <= 5'b01011; end
				10'b1011100011: begin sigmoid <= 7'b0001100; sigmoid_prime <= 5'b01011; end
				10'b1011100100: begin sigmoid <= 7'b0001101; sigmoid_prime <= 5'b01011; end
				10'b1011100101: begin sigmoid <= 7'b0001101; sigmoid_prime <= 5'b01011; end
				10'b1011100110: begin sigmoid <= 7'b0001101; sigmoid_prime <= 5'b01011; end
				10'b1011100111: begin sigmoid <= 7'b0001101; sigmoid_prime <= 5'b01100; end
				10'b1011101000: begin sigmoid <= 7'b0001101; sigmoid_prime <= 5'b01100; end
				10'b1011101001: begin sigmoid <= 7'b0001101; sigmoid_prime <= 5'b01100; end
				10'b1011101010: begin sigmoid <= 7'b0001101; sigmoid_prime <= 5'b01100; end
				10'b1011101011: begin sigmoid <= 7'b0001101; sigmoid_prime <= 5'b01100; end
				10'b1011101100: begin sigmoid <= 7'b0001101; sigmoid_prime <= 5'b01100; end
				10'b1011101101: begin sigmoid <= 7'b0001101; sigmoid_prime <= 5'b01100; end
				10'b1011101110: begin sigmoid <= 7'b0001101; sigmoid_prime <= 5'b01100; end
				10'b1011101111: begin sigmoid <= 7'b0001110; sigmoid_prime <= 5'b01100; end
				10'b1011110000: begin sigmoid <= 7'b0001110; sigmoid_prime <= 5'b01100; end
				10'b1011110001: begin sigmoid <= 7'b0001110; sigmoid_prime <= 5'b01100; end
				10'b1011110010: begin sigmoid <= 7'b0001110; sigmoid_prime <= 5'b01100; end
				10'b1011110011: begin sigmoid <= 7'b0001110; sigmoid_prime <= 5'b01100; end
				10'b1011110100: begin sigmoid <= 7'b0001110; sigmoid_prime <= 5'b01101; end
				10'b1011110101: begin sigmoid <= 7'b0001110; sigmoid_prime <= 5'b01101; end
				10'b1011110110: begin sigmoid <= 7'b0001110; sigmoid_prime <= 5'b01101; end
				10'b1011110111: begin sigmoid <= 7'b0001110; sigmoid_prime <= 5'b01101; end
				10'b1011111000: begin sigmoid <= 7'b0001110; sigmoid_prime <= 5'b01101; end
				10'b1011111001: begin sigmoid <= 7'b0001111; sigmoid_prime <= 5'b01101; end
				10'b1011111010: begin sigmoid <= 7'b0001111; sigmoid_prime <= 5'b01101; end
				10'b1011111011: begin sigmoid <= 7'b0001111; sigmoid_prime <= 5'b01101; end
				10'b1011111100: begin sigmoid <= 7'b0001111; sigmoid_prime <= 5'b01101; end
				10'b1011111101: begin sigmoid <= 7'b0001111; sigmoid_prime <= 5'b01101; end
				10'b1011111110: begin sigmoid <= 7'b0001111; sigmoid_prime <= 5'b01101; end
				10'b1011111111: begin sigmoid <= 7'b0001111; sigmoid_prime <= 5'b01101; end
				10'b1100000000: begin sigmoid <= 7'b0001111; sigmoid_prime <= 5'b01101; end
				10'b1100000001: begin sigmoid <= 7'b0001111; sigmoid_prime <= 5'b01110; end
				10'b1100000010: begin sigmoid <= 7'b0001111; sigmoid_prime <= 5'b01110; end
				10'b1100000011: begin sigmoid <= 7'b0010000; sigmoid_prime <= 5'b01110; end
				10'b1100000100: begin sigmoid <= 7'b0010000; sigmoid_prime <= 5'b01110; end
				10'b1100000101: begin sigmoid <= 7'b0010000; sigmoid_prime <= 5'b01110; end
				10'b1100000110: begin sigmoid <= 7'b0010000; sigmoid_prime <= 5'b01110; end
				10'b1100000111: begin sigmoid <= 7'b0010000; sigmoid_prime <= 5'b01110; end
				10'b1100001000: begin sigmoid <= 7'b0010000; sigmoid_prime <= 5'b01110; end
				10'b1100001001: begin sigmoid <= 7'b0010000; sigmoid_prime <= 5'b01110; end
				10'b1100001010: begin sigmoid <= 7'b0010000; sigmoid_prime <= 5'b01110; end
				10'b1100001011: begin sigmoid <= 7'b0010000; sigmoid_prime <= 5'b01110; end
				10'b1100001100: begin sigmoid <= 7'b0010001; sigmoid_prime <= 5'b01110; end
				10'b1100001101: begin sigmoid <= 7'b0010001; sigmoid_prime <= 5'b01111; end
				10'b1100001110: begin sigmoid <= 7'b0010001; sigmoid_prime <= 5'b01111; end
				10'b1100001111: begin sigmoid <= 7'b0010001; sigmoid_prime <= 5'b01111; end
				10'b1100010000: begin sigmoid <= 7'b0010001; sigmoid_prime <= 5'b01111; end
				10'b1100010001: begin sigmoid <= 7'b0010001; sigmoid_prime <= 5'b01111; end
				10'b1100010010: begin sigmoid <= 7'b0010001; sigmoid_prime <= 5'b01111; end
				10'b1100010011: begin sigmoid <= 7'b0010001; sigmoid_prime <= 5'b01111; end
				10'b1100010100: begin sigmoid <= 7'b0010001; sigmoid_prime <= 5'b01111; end
				10'b1100010101: begin sigmoid <= 7'b0010010; sigmoid_prime <= 5'b01111; end
				10'b1100010110: begin sigmoid <= 7'b0010010; sigmoid_prime <= 5'b01111; end
				10'b1100010111: begin sigmoid <= 7'b0010010; sigmoid_prime <= 5'b01111; end
				10'b1100011000: begin sigmoid <= 7'b0010010; sigmoid_prime <= 5'b01111; end
				10'b1100011001: begin sigmoid <= 7'b0010010; sigmoid_prime <= 5'b10000; end
				10'b1100011010: begin sigmoid <= 7'b0010010; sigmoid_prime <= 5'b10000; end
				10'b1100011011: begin sigmoid <= 7'b0010010; sigmoid_prime <= 5'b10000; end
				10'b1100011100: begin sigmoid <= 7'b0010010; sigmoid_prime <= 5'b10000; end
				10'b1100011101: begin sigmoid <= 7'b0010011; sigmoid_prime <= 5'b10000; end
				10'b1100011110: begin sigmoid <= 7'b0010011; sigmoid_prime <= 5'b10000; end
				10'b1100011111: begin sigmoid <= 7'b0010011; sigmoid_prime <= 5'b10000; end
				10'b1100100000: begin sigmoid <= 7'b0010011; sigmoid_prime <= 5'b10000; end
				10'b1100100001: begin sigmoid <= 7'b0010011; sigmoid_prime <= 5'b10000; end
				10'b1100100010: begin sigmoid <= 7'b0010011; sigmoid_prime <= 5'b10000; end
				10'b1100100011: begin sigmoid <= 7'b0010011; sigmoid_prime <= 5'b10000; end
				10'b1100100100: begin sigmoid <= 7'b0010011; sigmoid_prime <= 5'b10001; end
				10'b1100100101: begin sigmoid <= 7'b0010100; sigmoid_prime <= 5'b10001; end
				10'b1100100110: begin sigmoid <= 7'b0010100; sigmoid_prime <= 5'b10001; end
				10'b1100100111: begin sigmoid <= 7'b0010100; sigmoid_prime <= 5'b10001; end
				10'b1100101000: begin sigmoid <= 7'b0010100; sigmoid_prime <= 5'b10001; end
				10'b1100101001: begin sigmoid <= 7'b0010100; sigmoid_prime <= 5'b10001; end
				10'b1100101010: begin sigmoid <= 7'b0010100; sigmoid_prime <= 5'b10001; end
				10'b1100101011: begin sigmoid <= 7'b0010100; sigmoid_prime <= 5'b10001; end
				10'b1100101100: begin sigmoid <= 7'b0010101; sigmoid_prime <= 5'b10001; end
				10'b1100101101: begin sigmoid <= 7'b0010101; sigmoid_prime <= 5'b10001; end
				10'b1100101110: begin sigmoid <= 7'b0010101; sigmoid_prime <= 5'b10001; end
				10'b1100101111: begin sigmoid <= 7'b0010101; sigmoid_prime <= 5'b10010; end
				10'b1100110000: begin sigmoid <= 7'b0010101; sigmoid_prime <= 5'b10010; end
				10'b1100110001: begin sigmoid <= 7'b0010101; sigmoid_prime <= 5'b10010; end
				10'b1100110010: begin sigmoid <= 7'b0010101; sigmoid_prime <= 5'b10010; end
				10'b1100110011: begin sigmoid <= 7'b0010101; sigmoid_prime <= 5'b10010; end
				10'b1100110100: begin sigmoid <= 7'b0010110; sigmoid_prime <= 5'b10010; end
				10'b1100110101: begin sigmoid <= 7'b0010110; sigmoid_prime <= 5'b10010; end
				10'b1100110110: begin sigmoid <= 7'b0010110; sigmoid_prime <= 5'b10010; end
				10'b1100110111: begin sigmoid <= 7'b0010110; sigmoid_prime <= 5'b10010; end
				10'b1100111000: begin sigmoid <= 7'b0010110; sigmoid_prime <= 5'b10010; end
				10'b1100111001: begin sigmoid <= 7'b0010110; sigmoid_prime <= 5'b10010; end
				10'b1100111010: begin sigmoid <= 7'b0010110; sigmoid_prime <= 5'b10011; end
				10'b1100111011: begin sigmoid <= 7'b0010111; sigmoid_prime <= 5'b10011; end
				10'b1100111100: begin sigmoid <= 7'b0010111; sigmoid_prime <= 5'b10011; end
				10'b1100111101: begin sigmoid <= 7'b0010111; sigmoid_prime <= 5'b10011; end
				10'b1100111110: begin sigmoid <= 7'b0010111; sigmoid_prime <= 5'b10011; end
				10'b1100111111: begin sigmoid <= 7'b0010111; sigmoid_prime <= 5'b10011; end
				10'b1101000000: begin sigmoid <= 7'b0010111; sigmoid_prime <= 5'b10011; end
				10'b1101000001: begin sigmoid <= 7'b0010111; sigmoid_prime <= 5'b10011; end
				10'b1101000010: begin sigmoid <= 7'b0011000; sigmoid_prime <= 5'b10011; end
				10'b1101000011: begin sigmoid <= 7'b0011000; sigmoid_prime <= 5'b10011; end
				10'b1101000100: begin sigmoid <= 7'b0011000; sigmoid_prime <= 5'b10011; end
				10'b1101000101: begin sigmoid <= 7'b0011000; sigmoid_prime <= 5'b10100; end
				10'b1101000110: begin sigmoid <= 7'b0011000; sigmoid_prime <= 5'b10100; end
				10'b1101000111: begin sigmoid <= 7'b0011000; sigmoid_prime <= 5'b10100; end
				10'b1101001000: begin sigmoid <= 7'b0011001; sigmoid_prime <= 5'b10100; end
				10'b1101001001: begin sigmoid <= 7'b0011001; sigmoid_prime <= 5'b10100; end
				10'b1101001010: begin sigmoid <= 7'b0011001; sigmoid_prime <= 5'b10100; end
				10'b1101001011: begin sigmoid <= 7'b0011001; sigmoid_prime <= 5'b10100; end
				10'b1101001100: begin sigmoid <= 7'b0011001; sigmoid_prime <= 5'b10100; end
				10'b1101001101: begin sigmoid <= 7'b0011001; sigmoid_prime <= 5'b10100; end
				10'b1101001110: begin sigmoid <= 7'b0011010; sigmoid_prime <= 5'b10100; end
				10'b1101001111: begin sigmoid <= 7'b0011010; sigmoid_prime <= 5'b10101; end
				10'b1101010000: begin sigmoid <= 7'b0011010; sigmoid_prime <= 5'b10101; end
				10'b1101010001: begin sigmoid <= 7'b0011010; sigmoid_prime <= 5'b10101; end
				10'b1101010010: begin sigmoid <= 7'b0011010; sigmoid_prime <= 5'b10101; end
				10'b1101010011: begin sigmoid <= 7'b0011010; sigmoid_prime <= 5'b10101; end
				10'b1101010100: begin sigmoid <= 7'b0011010; sigmoid_prime <= 5'b10101; end
				10'b1101010101: begin sigmoid <= 7'b0011011; sigmoid_prime <= 5'b10101; end
				10'b1101010110: begin sigmoid <= 7'b0011011; sigmoid_prime <= 5'b10101; end
				10'b1101010111: begin sigmoid <= 7'b0011011; sigmoid_prime <= 5'b10101; end
				10'b1101011000: begin sigmoid <= 7'b0011011; sigmoid_prime <= 5'b10101; end
				10'b1101011001: begin sigmoid <= 7'b0011011; sigmoid_prime <= 5'b10101; end
				10'b1101011010: begin sigmoid <= 7'b0011011; sigmoid_prime <= 5'b10110; end
				10'b1101011011: begin sigmoid <= 7'b0011100; sigmoid_prime <= 5'b10110; end
				10'b1101011100: begin sigmoid <= 7'b0011100; sigmoid_prime <= 5'b10110; end
				10'b1101011101: begin sigmoid <= 7'b0011100; sigmoid_prime <= 5'b10110; end
				10'b1101011110: begin sigmoid <= 7'b0011100; sigmoid_prime <= 5'b10110; end
				10'b1101011111: begin sigmoid <= 7'b0011100; sigmoid_prime <= 5'b10110; end
				10'b1101100000: begin sigmoid <= 7'b0011101; sigmoid_prime <= 5'b10110; end
				10'b1101100001: begin sigmoid <= 7'b0011101; sigmoid_prime <= 5'b10110; end
				10'b1101100010: begin sigmoid <= 7'b0011101; sigmoid_prime <= 5'b10110; end
				10'b1101100011: begin sigmoid <= 7'b0011101; sigmoid_prime <= 5'b10110; end
				10'b1101100100: begin sigmoid <= 7'b0011101; sigmoid_prime <= 5'b10111; end
				10'b1101100101: begin sigmoid <= 7'b0011101; sigmoid_prime <= 5'b10111; end
				10'b1101100110: begin sigmoid <= 7'b0011110; sigmoid_prime <= 5'b10111; end
				10'b1101100111: begin sigmoid <= 7'b0011110; sigmoid_prime <= 5'b10111; end
				10'b1101101000: begin sigmoid <= 7'b0011110; sigmoid_prime <= 5'b10111; end
				10'b1101101001: begin sigmoid <= 7'b0011110; sigmoid_prime <= 5'b10111; end
				10'b1101101010: begin sigmoid <= 7'b0011110; sigmoid_prime <= 5'b10111; end
				10'b1101101011: begin sigmoid <= 7'b0011110; sigmoid_prime <= 5'b10111; end
				10'b1101101100: begin sigmoid <= 7'b0011111; sigmoid_prime <= 5'b10111; end
				10'b1101101101: begin sigmoid <= 7'b0011111; sigmoid_prime <= 5'b10111; end
				10'b1101101110: begin sigmoid <= 7'b0011111; sigmoid_prime <= 5'b10111; end
				10'b1101101111: begin sigmoid <= 7'b0011111; sigmoid_prime <= 5'b11000; end
				10'b1101110000: begin sigmoid <= 7'b0011111; sigmoid_prime <= 5'b11000; end
				10'b1101110001: begin sigmoid <= 7'b0100000; sigmoid_prime <= 5'b11000; end
				10'b1101110010: begin sigmoid <= 7'b0100000; sigmoid_prime <= 5'b11000; end
				10'b1101110011: begin sigmoid <= 7'b0100000; sigmoid_prime <= 5'b11000; end
				10'b1101110100: begin sigmoid <= 7'b0100000; sigmoid_prime <= 5'b11000; end
				10'b1101110101: begin sigmoid <= 7'b0100000; sigmoid_prime <= 5'b11000; end
				10'b1101110110: begin sigmoid <= 7'b0100000; sigmoid_prime <= 5'b11000; end
				10'b1101110111: begin sigmoid <= 7'b0100001; sigmoid_prime <= 5'b11000; end
				10'b1101111000: begin sigmoid <= 7'b0100001; sigmoid_prime <= 5'b11000; end
				10'b1101111001: begin sigmoid <= 7'b0100001; sigmoid_prime <= 5'b11001; end
				10'b1101111010: begin sigmoid <= 7'b0100001; sigmoid_prime <= 5'b11001; end
				10'b1101111011: begin sigmoid <= 7'b0100001; sigmoid_prime <= 5'b11001; end
				10'b1101111100: begin sigmoid <= 7'b0100010; sigmoid_prime <= 5'b11001; end
				10'b1101111101: begin sigmoid <= 7'b0100010; sigmoid_prime <= 5'b11001; end
				10'b1101111110: begin sigmoid <= 7'b0100010; sigmoid_prime <= 5'b11001; end
				10'b1101111111: begin sigmoid <= 7'b0100010; sigmoid_prime <= 5'b11001; end
				10'b1110000000: begin sigmoid <= 7'b0100010; sigmoid_prime <= 5'b11001; end
				10'b1110000001: begin sigmoid <= 7'b0100011; sigmoid_prime <= 5'b11001; end
				10'b1110000010: begin sigmoid <= 7'b0100011; sigmoid_prime <= 5'b11001; end
				10'b1110000011: begin sigmoid <= 7'b0100011; sigmoid_prime <= 5'b11001; end
				10'b1110000100: begin sigmoid <= 7'b0100011; sigmoid_prime <= 5'b11010; end
				10'b1110000101: begin sigmoid <= 7'b0100011; sigmoid_prime <= 5'b11010; end
				10'b1110000110: begin sigmoid <= 7'b0100100; sigmoid_prime <= 5'b11010; end
				10'b1110000111: begin sigmoid <= 7'b0100100; sigmoid_prime <= 5'b11010; end
				10'b1110001000: begin sigmoid <= 7'b0100100; sigmoid_prime <= 5'b11010; end
				10'b1110001001: begin sigmoid <= 7'b0100100; sigmoid_prime <= 5'b11010; end
				10'b1110001010: begin sigmoid <= 7'b0100100; sigmoid_prime <= 5'b11010; end
				10'b1110001011: begin sigmoid <= 7'b0100101; sigmoid_prime <= 5'b11010; end
				10'b1110001100: begin sigmoid <= 7'b0100101; sigmoid_prime <= 5'b11010; end
				10'b1110001101: begin sigmoid <= 7'b0100101; sigmoid_prime <= 5'b11010; end
				10'b1110001110: begin sigmoid <= 7'b0100101; sigmoid_prime <= 5'b11010; end
				10'b1110001111: begin sigmoid <= 7'b0100101; sigmoid_prime <= 5'b11010; end
				10'b1110010000: begin sigmoid <= 7'b0100110; sigmoid_prime <= 5'b11011; end
				10'b1110010001: begin sigmoid <= 7'b0100110; sigmoid_prime <= 5'b11011; end
				10'b1110010010: begin sigmoid <= 7'b0100110; sigmoid_prime <= 5'b11011; end
				10'b1110010011: begin sigmoid <= 7'b0100110; sigmoid_prime <= 5'b11011; end
				10'b1110010100: begin sigmoid <= 7'b0100110; sigmoid_prime <= 5'b11011; end
				10'b1110010101: begin sigmoid <= 7'b0100111; sigmoid_prime <= 5'b11011; end
				10'b1110010110: begin sigmoid <= 7'b0100111; sigmoid_prime <= 5'b11011; end
				10'b1110010111: begin sigmoid <= 7'b0100111; sigmoid_prime <= 5'b11011; end
				10'b1110011000: begin sigmoid <= 7'b0100111; sigmoid_prime <= 5'b11011; end
				10'b1110011001: begin sigmoid <= 7'b0101000; sigmoid_prime <= 5'b11011; end
				10'b1110011010: begin sigmoid <= 7'b0101000; sigmoid_prime <= 5'b11011; end
				10'b1110011011: begin sigmoid <= 7'b0101000; sigmoid_prime <= 5'b11011; end
				10'b1110011100: begin sigmoid <= 7'b0101000; sigmoid_prime <= 5'b11100; end
				10'b1110011101: begin sigmoid <= 7'b0101000; sigmoid_prime <= 5'b11100; end
				10'b1110011110: begin sigmoid <= 7'b0101001; sigmoid_prime <= 5'b11100; end
				10'b1110011111: begin sigmoid <= 7'b0101001; sigmoid_prime <= 5'b11100; end
				10'b1110100000: begin sigmoid <= 7'b0101001; sigmoid_prime <= 5'b11100; end
				10'b1110100001: begin sigmoid <= 7'b0101001; sigmoid_prime <= 5'b11100; end
				10'b1110100010: begin sigmoid <= 7'b0101010; sigmoid_prime <= 5'b11100; end
				10'b1110100011: begin sigmoid <= 7'b0101010; sigmoid_prime <= 5'b11100; end
				10'b1110100100: begin sigmoid <= 7'b0101010; sigmoid_prime <= 5'b11100; end
				10'b1110100101: begin sigmoid <= 7'b0101010; sigmoid_prime <= 5'b11100; end
				10'b1110100110: begin sigmoid <= 7'b0101010; sigmoid_prime <= 5'b11100; end
				10'b1110100111: begin sigmoid <= 7'b0101011; sigmoid_prime <= 5'b11100; end
				10'b1110101000: begin sigmoid <= 7'b0101011; sigmoid_prime <= 5'b11100; end
				10'b1110101001: begin sigmoid <= 7'b0101011; sigmoid_prime <= 5'b11101; end
				10'b1110101010: begin sigmoid <= 7'b0101011; sigmoid_prime <= 5'b11101; end
				10'b1110101011: begin sigmoid <= 7'b0101011; sigmoid_prime <= 5'b11101; end
				10'b1110101100: begin sigmoid <= 7'b0101100; sigmoid_prime <= 5'b11101; end
				10'b1110101101: begin sigmoid <= 7'b0101100; sigmoid_prime <= 5'b11101; end
				10'b1110101110: begin sigmoid <= 7'b0101100; sigmoid_prime <= 5'b11101; end
				10'b1110101111: begin sigmoid <= 7'b0101100; sigmoid_prime <= 5'b11101; end
				10'b1110110000: begin sigmoid <= 7'b0101101; sigmoid_prime <= 5'b11101; end
				10'b1110110001: begin sigmoid <= 7'b0101101; sigmoid_prime <= 5'b11101; end
				10'b1110110010: begin sigmoid <= 7'b0101101; sigmoid_prime <= 5'b11101; end
				10'b1110110011: begin sigmoid <= 7'b0101101; sigmoid_prime <= 5'b11101; end
				10'b1110110100: begin sigmoid <= 7'b0101110; sigmoid_prime <= 5'b11101; end
				10'b1110110101: begin sigmoid <= 7'b0101110; sigmoid_prime <= 5'b11101; end
				10'b1110110110: begin sigmoid <= 7'b0101110; sigmoid_prime <= 5'b11101; end
				10'b1110110111: begin sigmoid <= 7'b0101110; sigmoid_prime <= 5'b11110; end
				10'b1110111000: begin sigmoid <= 7'b0101110; sigmoid_prime <= 5'b11110; end
				10'b1110111001: begin sigmoid <= 7'b0101111; sigmoid_prime <= 5'b11110; end
				10'b1110111010: begin sigmoid <= 7'b0101111; sigmoid_prime <= 5'b11110; end
				10'b1110111011: begin sigmoid <= 7'b0101111; sigmoid_prime <= 5'b11110; end
				10'b1110111100: begin sigmoid <= 7'b0101111; sigmoid_prime <= 5'b11110; end
				10'b1110111101: begin sigmoid <= 7'b0110000; sigmoid_prime <= 5'b11110; end
				10'b1110111110: begin sigmoid <= 7'b0110000; sigmoid_prime <= 5'b11110; end
				10'b1110111111: begin sigmoid <= 7'b0110000; sigmoid_prime <= 5'b11110; end
				10'b1111000000: begin sigmoid <= 7'b0110000; sigmoid_prime <= 5'b11110; end
				10'b1111000001: begin sigmoid <= 7'b0110001; sigmoid_prime <= 5'b11110; end
				10'b1111000010: begin sigmoid <= 7'b0110001; sigmoid_prime <= 5'b11110; end
				10'b1111000011: begin sigmoid <= 7'b0110001; sigmoid_prime <= 5'b11110; end
				10'b1111000100: begin sigmoid <= 7'b0110001; sigmoid_prime <= 5'b11110; end
				10'b1111000101: begin sigmoid <= 7'b0110010; sigmoid_prime <= 5'b11110; end
				10'b1111000110: begin sigmoid <= 7'b0110010; sigmoid_prime <= 5'b11110; end
				10'b1111000111: begin sigmoid <= 7'b0110010; sigmoid_prime <= 5'b11110; end
				10'b1111001000: begin sigmoid <= 7'b0110010; sigmoid_prime <= 5'b11111; end
				10'b1111001001: begin sigmoid <= 7'b0110010; sigmoid_prime <= 5'b11111; end
				10'b1111001010: begin sigmoid <= 7'b0110011; sigmoid_prime <= 5'b11111; end
				10'b1111001011: begin sigmoid <= 7'b0110011; sigmoid_prime <= 5'b11111; end
				10'b1111001100: begin sigmoid <= 7'b0110011; sigmoid_prime <= 5'b11111; end
				10'b1111001101: begin sigmoid <= 7'b0110011; sigmoid_prime <= 5'b11111; end
				10'b1111001110: begin sigmoid <= 7'b0110100; sigmoid_prime <= 5'b11111; end
				10'b1111001111: begin sigmoid <= 7'b0110100; sigmoid_prime <= 5'b11111; end
				10'b1111010000: begin sigmoid <= 7'b0110100; sigmoid_prime <= 5'b11111; end
				10'b1111010001: begin sigmoid <= 7'b0110100; sigmoid_prime <= 5'b11111; end
				10'b1111010010: begin sigmoid <= 7'b0110101; sigmoid_prime <= 5'b11111; end
				10'b1111010011: begin sigmoid <= 7'b0110101; sigmoid_prime <= 5'b11111; end
				10'b1111010100: begin sigmoid <= 7'b0110101; sigmoid_prime <= 5'b11111; end
				10'b1111010101: begin sigmoid <= 7'b0110101; sigmoid_prime <= 5'b11111; end
				10'b1111010110: begin sigmoid <= 7'b0110110; sigmoid_prime <= 5'b11111; end
				10'b1111010111: begin sigmoid <= 7'b0110110; sigmoid_prime <= 5'b11111; end
				10'b1111011000: begin sigmoid <= 7'b0110110; sigmoid_prime <= 5'b11111; end
				10'b1111011001: begin sigmoid <= 7'b0110110; sigmoid_prime <= 5'b11111; end
				10'b1111011010: begin sigmoid <= 7'b0110111; sigmoid_prime <= 5'b11111; end
				10'b1111011011: begin sigmoid <= 7'b0110111; sigmoid_prime <= 5'b11111; end
				10'b1111011100: begin sigmoid <= 7'b0110111; sigmoid_prime <= 5'b11111; end
				10'b1111011101: begin sigmoid <= 7'b0110111; sigmoid_prime <= 5'b11111; end
				10'b1111011110: begin sigmoid <= 7'b0111000; sigmoid_prime <= 5'b11111; end
				10'b1111011111: begin sigmoid <= 7'b0111000; sigmoid_prime <= 5'b11111; end
				10'b1111100000: begin sigmoid <= 7'b0111000; sigmoid_prime <= 5'b11111; end
				10'b1111100001: begin sigmoid <= 7'b0111000; sigmoid_prime <= 5'b11111; end
				10'b1111100010: begin sigmoid <= 7'b0111001; sigmoid_prime <= 5'b11111; end
				10'b1111100011: begin sigmoid <= 7'b0111001; sigmoid_prime <= 5'b11111; end
				10'b1111100100: begin sigmoid <= 7'b0111001; sigmoid_prime <= 5'b11111; end
				10'b1111100101: begin sigmoid <= 7'b0111001; sigmoid_prime <= 5'b11111; end
				10'b1111100110: begin sigmoid <= 7'b0111010; sigmoid_prime <= 5'b11111; end
				10'b1111100111: begin sigmoid <= 7'b0111010; sigmoid_prime <= 5'b11111; end
				10'b1111101000: begin sigmoid <= 7'b0111010; sigmoid_prime <= 5'b11111; end
				10'b1111101001: begin sigmoid <= 7'b0111010; sigmoid_prime <= 5'b11111; end
				10'b1111101010: begin sigmoid <= 7'b0111011; sigmoid_prime <= 5'b11111; end
				10'b1111101011: begin sigmoid <= 7'b0111011; sigmoid_prime <= 5'b11111; end
				10'b1111101100: begin sigmoid <= 7'b0111011; sigmoid_prime <= 5'b11111; end
				10'b1111101101: begin sigmoid <= 7'b0111011; sigmoid_prime <= 5'b11111; end
				10'b1111101110: begin sigmoid <= 7'b0111100; sigmoid_prime <= 5'b11111; end
				10'b1111101111: begin sigmoid <= 7'b0111100; sigmoid_prime <= 5'b11111; end
				10'b1111110000: begin sigmoid <= 7'b0111100; sigmoid_prime <= 5'b11111; end
				10'b1111110001: begin sigmoid <= 7'b0111100; sigmoid_prime <= 5'b11111; end
				10'b1111110010: begin sigmoid <= 7'b0111101; sigmoid_prime <= 5'b11111; end
				10'b1111110011: begin sigmoid <= 7'b0111101; sigmoid_prime <= 5'b11111; end
				10'b1111110100: begin sigmoid <= 7'b0111101; sigmoid_prime <= 5'b11111; end
				10'b1111110101: begin sigmoid <= 7'b0111101; sigmoid_prime <= 5'b11111; end
				10'b1111110110: begin sigmoid <= 7'b0111110; sigmoid_prime <= 5'b11111; end
				10'b1111110111: begin sigmoid <= 7'b0111110; sigmoid_prime <= 5'b11111; end
				10'b1111111000: begin sigmoid <= 7'b0111110; sigmoid_prime <= 5'b11111; end
				10'b1111111001: begin sigmoid <= 7'b0111110; sigmoid_prime <= 5'b11111; end
				10'b1111111010: begin sigmoid <= 7'b0111111; sigmoid_prime <= 5'b11111; end
				10'b1111111011: begin sigmoid <= 7'b0111111; sigmoid_prime <= 5'b11111; end
				10'b1111111100: begin sigmoid <= 7'b0111111; sigmoid_prime <= 5'b11111; end
				10'b1111111101: begin sigmoid <= 7'b0111111; sigmoid_prime <= 5'b11111; end
				10'b1111111110: begin sigmoid <= 7'b1000000; sigmoid_prime <= 5'b11111; end
				10'b1111111111: begin sigmoid <= 7'b1000000; sigmoid_prime <= 5'b11111; end
				10'b0000000000: begin sigmoid <= 7'b1000000; sigmoid_prime <= 5'b11111; end
				10'b0000000001: begin sigmoid <= 7'b1000000; sigmoid_prime <= 5'b11111; end
				10'b0000000010: begin sigmoid <= 7'b1000000; sigmoid_prime <= 5'b11111; end
				10'b0000000011: begin sigmoid <= 7'b1000001; sigmoid_prime <= 5'b11111; end
				10'b0000000100: begin sigmoid <= 7'b1000001; sigmoid_prime <= 5'b11111; end
				10'b0000000101: begin sigmoid <= 7'b1000001; sigmoid_prime <= 5'b11111; end
				10'b0000000110: begin sigmoid <= 7'b1000001; sigmoid_prime <= 5'b11111; end
				10'b0000000111: begin sigmoid <= 7'b1000010; sigmoid_prime <= 5'b11111; end
				10'b0000001000: begin sigmoid <= 7'b1000010; sigmoid_prime <= 5'b11111; end
				10'b0000001001: begin sigmoid <= 7'b1000010; sigmoid_prime <= 5'b11111; end
				10'b0000001010: begin sigmoid <= 7'b1000010; sigmoid_prime <= 5'b11111; end
				10'b0000001011: begin sigmoid <= 7'b1000011; sigmoid_prime <= 5'b11111; end
				10'b0000001100: begin sigmoid <= 7'b1000011; sigmoid_prime <= 5'b11111; end
				10'b0000001101: begin sigmoid <= 7'b1000011; sigmoid_prime <= 5'b11111; end
				10'b0000001110: begin sigmoid <= 7'b1000011; sigmoid_prime <= 5'b11111; end
				10'b0000001111: begin sigmoid <= 7'b1000100; sigmoid_prime <= 5'b11111; end
				10'b0000010000: begin sigmoid <= 7'b1000100; sigmoid_prime <= 5'b11111; end
				10'b0000010001: begin sigmoid <= 7'b1000100; sigmoid_prime <= 5'b11111; end
				10'b0000010010: begin sigmoid <= 7'b1000100; sigmoid_prime <= 5'b11111; end
				10'b0000010011: begin sigmoid <= 7'b1000101; sigmoid_prime <= 5'b11111; end
				10'b0000010100: begin sigmoid <= 7'b1000101; sigmoid_prime <= 5'b11111; end
				10'b0000010101: begin sigmoid <= 7'b1000101; sigmoid_prime <= 5'b11111; end
				10'b0000010110: begin sigmoid <= 7'b1000101; sigmoid_prime <= 5'b11111; end
				10'b0000010111: begin sigmoid <= 7'b1000110; sigmoid_prime <= 5'b11111; end
				10'b0000011000: begin sigmoid <= 7'b1000110; sigmoid_prime <= 5'b11111; end
				10'b0000011001: begin sigmoid <= 7'b1000110; sigmoid_prime <= 5'b11111; end
				10'b0000011010: begin sigmoid <= 7'b1000110; sigmoid_prime <= 5'b11111; end
				10'b0000011011: begin sigmoid <= 7'b1000111; sigmoid_prime <= 5'b11111; end
				10'b0000011100: begin sigmoid <= 7'b1000111; sigmoid_prime <= 5'b11111; end
				10'b0000011101: begin sigmoid <= 7'b1000111; sigmoid_prime <= 5'b11111; end
				10'b0000011110: begin sigmoid <= 7'b1000111; sigmoid_prime <= 5'b11111; end
				10'b0000011111: begin sigmoid <= 7'b1001000; sigmoid_prime <= 5'b11111; end
				10'b0000100000: begin sigmoid <= 7'b1001000; sigmoid_prime <= 5'b11111; end
				10'b0000100001: begin sigmoid <= 7'b1001000; sigmoid_prime <= 5'b11111; end
				10'b0000100010: begin sigmoid <= 7'b1001000; sigmoid_prime <= 5'b11111; end
				10'b0000100011: begin sigmoid <= 7'b1001001; sigmoid_prime <= 5'b11111; end
				10'b0000100100: begin sigmoid <= 7'b1001001; sigmoid_prime <= 5'b11111; end
				10'b0000100101: begin sigmoid <= 7'b1001001; sigmoid_prime <= 5'b11111; end
				10'b0000100110: begin sigmoid <= 7'b1001001; sigmoid_prime <= 5'b11111; end
				10'b0000100111: begin sigmoid <= 7'b1001010; sigmoid_prime <= 5'b11111; end
				10'b0000101000: begin sigmoid <= 7'b1001010; sigmoid_prime <= 5'b11111; end
				10'b0000101001: begin sigmoid <= 7'b1001010; sigmoid_prime <= 5'b11111; end
				10'b0000101010: begin sigmoid <= 7'b1001010; sigmoid_prime <= 5'b11111; end
				10'b0000101011: begin sigmoid <= 7'b1001011; sigmoid_prime <= 5'b11111; end
				10'b0000101100: begin sigmoid <= 7'b1001011; sigmoid_prime <= 5'b11111; end
				10'b0000101101: begin sigmoid <= 7'b1001011; sigmoid_prime <= 5'b11111; end
				10'b0000101110: begin sigmoid <= 7'b1001011; sigmoid_prime <= 5'b11111; end
				10'b0000101111: begin sigmoid <= 7'b1001100; sigmoid_prime <= 5'b11111; end
				10'b0000110000: begin sigmoid <= 7'b1001100; sigmoid_prime <= 5'b11111; end
				10'b0000110001: begin sigmoid <= 7'b1001100; sigmoid_prime <= 5'b11111; end
				10'b0000110010: begin sigmoid <= 7'b1001100; sigmoid_prime <= 5'b11111; end
				10'b0000110011: begin sigmoid <= 7'b1001101; sigmoid_prime <= 5'b11111; end
				10'b0000110100: begin sigmoid <= 7'b1001101; sigmoid_prime <= 5'b11111; end
				10'b0000110101: begin sigmoid <= 7'b1001101; sigmoid_prime <= 5'b11111; end
				10'b0000110110: begin sigmoid <= 7'b1001101; sigmoid_prime <= 5'b11111; end
				10'b0000110111: begin sigmoid <= 7'b1001110; sigmoid_prime <= 5'b11111; end
				10'b0000111000: begin sigmoid <= 7'b1001110; sigmoid_prime <= 5'b11111; end
				10'b0000111001: begin sigmoid <= 7'b1001110; sigmoid_prime <= 5'b11110; end
				10'b0000111010: begin sigmoid <= 7'b1001110; sigmoid_prime <= 5'b11110; end
				10'b0000111011: begin sigmoid <= 7'b1001110; sigmoid_prime <= 5'b11110; end
				10'b0000111100: begin sigmoid <= 7'b1001111; sigmoid_prime <= 5'b11110; end
				10'b0000111101: begin sigmoid <= 7'b1001111; sigmoid_prime <= 5'b11110; end
				10'b0000111110: begin sigmoid <= 7'b1001111; sigmoid_prime <= 5'b11110; end
				10'b0000111111: begin sigmoid <= 7'b1001111; sigmoid_prime <= 5'b11110; end
				10'b0001000000: begin sigmoid <= 7'b1010000; sigmoid_prime <= 5'b11110; end
				10'b0001000001: begin sigmoid <= 7'b1010000; sigmoid_prime <= 5'b11110; end
				10'b0001000010: begin sigmoid <= 7'b1010000; sigmoid_prime <= 5'b11110; end
				10'b0001000011: begin sigmoid <= 7'b1010000; sigmoid_prime <= 5'b11110; end
				10'b0001000100: begin sigmoid <= 7'b1010001; sigmoid_prime <= 5'b11110; end
				10'b0001000101: begin sigmoid <= 7'b1010001; sigmoid_prime <= 5'b11110; end
				10'b0001000110: begin sigmoid <= 7'b1010001; sigmoid_prime <= 5'b11110; end
				10'b0001000111: begin sigmoid <= 7'b1010001; sigmoid_prime <= 5'b11110; end
				10'b0001001000: begin sigmoid <= 7'b1010010; sigmoid_prime <= 5'b11110; end
				10'b0001001001: begin sigmoid <= 7'b1010010; sigmoid_prime <= 5'b11110; end
				10'b0001001010: begin sigmoid <= 7'b1010010; sigmoid_prime <= 5'b11101; end
				10'b0001001011: begin sigmoid <= 7'b1010010; sigmoid_prime <= 5'b11101; end
				10'b0001001100: begin sigmoid <= 7'b1010010; sigmoid_prime <= 5'b11101; end
				10'b0001001101: begin sigmoid <= 7'b1010011; sigmoid_prime <= 5'b11101; end
				10'b0001001110: begin sigmoid <= 7'b1010011; sigmoid_prime <= 5'b11101; end
				10'b0001001111: begin sigmoid <= 7'b1010011; sigmoid_prime <= 5'b11101; end
				10'b0001010000: begin sigmoid <= 7'b1010011; sigmoid_prime <= 5'b11101; end
				10'b0001010001: begin sigmoid <= 7'b1010100; sigmoid_prime <= 5'b11101; end
				10'b0001010010: begin sigmoid <= 7'b1010100; sigmoid_prime <= 5'b11101; end
				10'b0001010011: begin sigmoid <= 7'b1010100; sigmoid_prime <= 5'b11101; end
				10'b0001010100: begin sigmoid <= 7'b1010100; sigmoid_prime <= 5'b11101; end
				10'b0001010101: begin sigmoid <= 7'b1010101; sigmoid_prime <= 5'b11101; end
				10'b0001010110: begin sigmoid <= 7'b1010101; sigmoid_prime <= 5'b11101; end
				10'b0001010111: begin sigmoid <= 7'b1010101; sigmoid_prime <= 5'b11101; end
				10'b0001011000: begin sigmoid <= 7'b1010101; sigmoid_prime <= 5'b11100; end
				10'b0001011001: begin sigmoid <= 7'b1010101; sigmoid_prime <= 5'b11100; end
				10'b0001011010: begin sigmoid <= 7'b1010110; sigmoid_prime <= 5'b11100; end
				10'b0001011011: begin sigmoid <= 7'b1010110; sigmoid_prime <= 5'b11100; end
				10'b0001011100: begin sigmoid <= 7'b1010110; sigmoid_prime <= 5'b11100; end
				10'b0001011101: begin sigmoid <= 7'b1010110; sigmoid_prime <= 5'b11100; end
				10'b0001011110: begin sigmoid <= 7'b1010110; sigmoid_prime <= 5'b11100; end
				10'b0001011111: begin sigmoid <= 7'b1010111; sigmoid_prime <= 5'b11100; end
				10'b0001100000: begin sigmoid <= 7'b1010111; sigmoid_prime <= 5'b11100; end
				10'b0001100001: begin sigmoid <= 7'b1010111; sigmoid_prime <= 5'b11100; end
				10'b0001100010: begin sigmoid <= 7'b1010111; sigmoid_prime <= 5'b11100; end
				10'b0001100011: begin sigmoid <= 7'b1011000; sigmoid_prime <= 5'b11100; end
				10'b0001100100: begin sigmoid <= 7'b1011000; sigmoid_prime <= 5'b11100; end
				10'b0001100101: begin sigmoid <= 7'b1011000; sigmoid_prime <= 5'b11011; end
				10'b0001100110: begin sigmoid <= 7'b1011000; sigmoid_prime <= 5'b11011; end
				10'b0001100111: begin sigmoid <= 7'b1011000; sigmoid_prime <= 5'b11011; end
				10'b0001101000: begin sigmoid <= 7'b1011001; sigmoid_prime <= 5'b11011; end
				10'b0001101001: begin sigmoid <= 7'b1011001; sigmoid_prime <= 5'b11011; end
				10'b0001101010: begin sigmoid <= 7'b1011001; sigmoid_prime <= 5'b11011; end
				10'b0001101011: begin sigmoid <= 7'b1011001; sigmoid_prime <= 5'b11011; end
				10'b0001101100: begin sigmoid <= 7'b1011010; sigmoid_prime <= 5'b11011; end
				10'b0001101101: begin sigmoid <= 7'b1011010; sigmoid_prime <= 5'b11011; end
				10'b0001101110: begin sigmoid <= 7'b1011010; sigmoid_prime <= 5'b11011; end
				10'b0001101111: begin sigmoid <= 7'b1011010; sigmoid_prime <= 5'b11011; end
				10'b0001110000: begin sigmoid <= 7'b1011010; sigmoid_prime <= 5'b11011; end
				10'b0001110001: begin sigmoid <= 7'b1011011; sigmoid_prime <= 5'b11010; end
				10'b0001110010: begin sigmoid <= 7'b1011011; sigmoid_prime <= 5'b11010; end
				10'b0001110011: begin sigmoid <= 7'b1011011; sigmoid_prime <= 5'b11010; end
				10'b0001110100: begin sigmoid <= 7'b1011011; sigmoid_prime <= 5'b11010; end
				10'b0001110101: begin sigmoid <= 7'b1011011; sigmoid_prime <= 5'b11010; end
				10'b0001110110: begin sigmoid <= 7'b1011100; sigmoid_prime <= 5'b11010; end
				10'b0001110111: begin sigmoid <= 7'b1011100; sigmoid_prime <= 5'b11010; end
				10'b0001111000: begin sigmoid <= 7'b1011100; sigmoid_prime <= 5'b11010; end
				10'b0001111001: begin sigmoid <= 7'b1011100; sigmoid_prime <= 5'b11010; end
				10'b0001111010: begin sigmoid <= 7'b1011100; sigmoid_prime <= 5'b11010; end
				10'b0001111011: begin sigmoid <= 7'b1011101; sigmoid_prime <= 5'b11010; end
				10'b0001111100: begin sigmoid <= 7'b1011101; sigmoid_prime <= 5'b11010; end
				10'b0001111101: begin sigmoid <= 7'b1011101; sigmoid_prime <= 5'b11001; end
				10'b0001111110: begin sigmoid <= 7'b1011101; sigmoid_prime <= 5'b11001; end
				10'b0001111111: begin sigmoid <= 7'b1011101; sigmoid_prime <= 5'b11001; end
				10'b0010000000: begin sigmoid <= 7'b1011110; sigmoid_prime <= 5'b11001; end
				10'b0010000001: begin sigmoid <= 7'b1011110; sigmoid_prime <= 5'b11001; end
				10'b0010000010: begin sigmoid <= 7'b1011110; sigmoid_prime <= 5'b11001; end
				10'b0010000011: begin sigmoid <= 7'b1011110; sigmoid_prime <= 5'b11001; end
				10'b0010000100: begin sigmoid <= 7'b1011110; sigmoid_prime <= 5'b11001; end
				10'b0010000101: begin sigmoid <= 7'b1011111; sigmoid_prime <= 5'b11001; end
				10'b0010000110: begin sigmoid <= 7'b1011111; sigmoid_prime <= 5'b11001; end
				10'b0010000111: begin sigmoid <= 7'b1011111; sigmoid_prime <= 5'b11001; end
				10'b0010001000: begin sigmoid <= 7'b1011111; sigmoid_prime <= 5'b11000; end
				10'b0010001001: begin sigmoid <= 7'b1011111; sigmoid_prime <= 5'b11000; end
				10'b0010001010: begin sigmoid <= 7'b1100000; sigmoid_prime <= 5'b11000; end
				10'b0010001011: begin sigmoid <= 7'b1100000; sigmoid_prime <= 5'b11000; end
				10'b0010001100: begin sigmoid <= 7'b1100000; sigmoid_prime <= 5'b11000; end
				10'b0010001101: begin sigmoid <= 7'b1100000; sigmoid_prime <= 5'b11000; end
				10'b0010001110: begin sigmoid <= 7'b1100000; sigmoid_prime <= 5'b11000; end
				10'b0010001111: begin sigmoid <= 7'b1100000; sigmoid_prime <= 5'b11000; end
				10'b0010010000: begin sigmoid <= 7'b1100001; sigmoid_prime <= 5'b11000; end
				10'b0010010001: begin sigmoid <= 7'b1100001; sigmoid_prime <= 5'b11000; end
				10'b0010010010: begin sigmoid <= 7'b1100001; sigmoid_prime <= 5'b10111; end
				10'b0010010011: begin sigmoid <= 7'b1100001; sigmoid_prime <= 5'b10111; end
				10'b0010010100: begin sigmoid <= 7'b1100001; sigmoid_prime <= 5'b10111; end
				10'b0010010101: begin sigmoid <= 7'b1100010; sigmoid_prime <= 5'b10111; end
				10'b0010010110: begin sigmoid <= 7'b1100010; sigmoid_prime <= 5'b10111; end
				10'b0010010111: begin sigmoid <= 7'b1100010; sigmoid_prime <= 5'b10111; end
				10'b0010011000: begin sigmoid <= 7'b1100010; sigmoid_prime <= 5'b10111; end
				10'b0010011001: begin sigmoid <= 7'b1100010; sigmoid_prime <= 5'b10111; end
				10'b0010011010: begin sigmoid <= 7'b1100010; sigmoid_prime <= 5'b10111; end
				10'b0010011011: begin sigmoid <= 7'b1100011; sigmoid_prime <= 5'b10111; end
				10'b0010011100: begin sigmoid <= 7'b1100011; sigmoid_prime <= 5'b10111; end
				10'b0010011101: begin sigmoid <= 7'b1100011; sigmoid_prime <= 5'b10110; end
				10'b0010011110: begin sigmoid <= 7'b1100011; sigmoid_prime <= 5'b10110; end
				10'b0010011111: begin sigmoid <= 7'b1100011; sigmoid_prime <= 5'b10110; end
				10'b0010100000: begin sigmoid <= 7'b1100011; sigmoid_prime <= 5'b10110; end
				10'b0010100001: begin sigmoid <= 7'b1100100; sigmoid_prime <= 5'b10110; end
				10'b0010100010: begin sigmoid <= 7'b1100100; sigmoid_prime <= 5'b10110; end
				10'b0010100011: begin sigmoid <= 7'b1100100; sigmoid_prime <= 5'b10110; end
				10'b0010100100: begin sigmoid <= 7'b1100100; sigmoid_prime <= 5'b10110; end
				10'b0010100101: begin sigmoid <= 7'b1100100; sigmoid_prime <= 5'b10110; end
				10'b0010100110: begin sigmoid <= 7'b1100101; sigmoid_prime <= 5'b10110; end
				10'b0010100111: begin sigmoid <= 7'b1100101; sigmoid_prime <= 5'b10101; end
				10'b0010101000: begin sigmoid <= 7'b1100101; sigmoid_prime <= 5'b10101; end
				10'b0010101001: begin sigmoid <= 7'b1100101; sigmoid_prime <= 5'b10101; end
				10'b0010101010: begin sigmoid <= 7'b1100101; sigmoid_prime <= 5'b10101; end
				10'b0010101011: begin sigmoid <= 7'b1100101; sigmoid_prime <= 5'b10101; end
				10'b0010101100: begin sigmoid <= 7'b1100110; sigmoid_prime <= 5'b10101; end
				10'b0010101101: begin sigmoid <= 7'b1100110; sigmoid_prime <= 5'b10101; end
				10'b0010101110: begin sigmoid <= 7'b1100110; sigmoid_prime <= 5'b10101; end
				10'b0010101111: begin sigmoid <= 7'b1100110; sigmoid_prime <= 5'b10101; end
				10'b0010110000: begin sigmoid <= 7'b1100110; sigmoid_prime <= 5'b10101; end
				10'b0010110001: begin sigmoid <= 7'b1100110; sigmoid_prime <= 5'b10101; end
				10'b0010110010: begin sigmoid <= 7'b1100110; sigmoid_prime <= 5'b10100; end
				10'b0010110011: begin sigmoid <= 7'b1100111; sigmoid_prime <= 5'b10100; end
				10'b0010110100: begin sigmoid <= 7'b1100111; sigmoid_prime <= 5'b10100; end
				10'b0010110101: begin sigmoid <= 7'b1100111; sigmoid_prime <= 5'b10100; end
				10'b0010110110: begin sigmoid <= 7'b1100111; sigmoid_prime <= 5'b10100; end
				10'b0010110111: begin sigmoid <= 7'b1100111; sigmoid_prime <= 5'b10100; end
				10'b0010111000: begin sigmoid <= 7'b1100111; sigmoid_prime <= 5'b10100; end
				10'b0010111001: begin sigmoid <= 7'b1101000; sigmoid_prime <= 5'b10100; end
				10'b0010111010: begin sigmoid <= 7'b1101000; sigmoid_prime <= 5'b10100; end
				10'b0010111011: begin sigmoid <= 7'b1101000; sigmoid_prime <= 5'b10100; end
				10'b0010111100: begin sigmoid <= 7'b1101000; sigmoid_prime <= 5'b10011; end
				10'b0010111101: begin sigmoid <= 7'b1101000; sigmoid_prime <= 5'b10011; end
				10'b0010111110: begin sigmoid <= 7'b1101000; sigmoid_prime <= 5'b10011; end
				10'b0010111111: begin sigmoid <= 7'b1101001; sigmoid_prime <= 5'b10011; end
				10'b0011000000: begin sigmoid <= 7'b1101001; sigmoid_prime <= 5'b10011; end
				10'b0011000001: begin sigmoid <= 7'b1101001; sigmoid_prime <= 5'b10011; end
				10'b0011000010: begin sigmoid <= 7'b1101001; sigmoid_prime <= 5'b10011; end
				10'b0011000011: begin sigmoid <= 7'b1101001; sigmoid_prime <= 5'b10011; end
				10'b0011000100: begin sigmoid <= 7'b1101001; sigmoid_prime <= 5'b10011; end
				10'b0011000101: begin sigmoid <= 7'b1101001; sigmoid_prime <= 5'b10011; end
				10'b0011000110: begin sigmoid <= 7'b1101010; sigmoid_prime <= 5'b10011; end
				10'b0011000111: begin sigmoid <= 7'b1101010; sigmoid_prime <= 5'b10010; end
				10'b0011001000: begin sigmoid <= 7'b1101010; sigmoid_prime <= 5'b10010; end
				10'b0011001001: begin sigmoid <= 7'b1101010; sigmoid_prime <= 5'b10010; end
				10'b0011001010: begin sigmoid <= 7'b1101010; sigmoid_prime <= 5'b10010; end
				10'b0011001011: begin sigmoid <= 7'b1101010; sigmoid_prime <= 5'b10010; end
				10'b0011001100: begin sigmoid <= 7'b1101010; sigmoid_prime <= 5'b10010; end
				10'b0011001101: begin sigmoid <= 7'b1101011; sigmoid_prime <= 5'b10010; end
				10'b0011001110: begin sigmoid <= 7'b1101011; sigmoid_prime <= 5'b10010; end
				10'b0011001111: begin sigmoid <= 7'b1101011; sigmoid_prime <= 5'b10010; end
				10'b0011010000: begin sigmoid <= 7'b1101011; sigmoid_prime <= 5'b10010; end
				10'b0011010001: begin sigmoid <= 7'b1101011; sigmoid_prime <= 5'b10010; end
				10'b0011010010: begin sigmoid <= 7'b1101011; sigmoid_prime <= 5'b10001; end
				10'b0011010011: begin sigmoid <= 7'b1101011; sigmoid_prime <= 5'b10001; end
				10'b0011010100: begin sigmoid <= 7'b1101011; sigmoid_prime <= 5'b10001; end
				10'b0011010101: begin sigmoid <= 7'b1101100; sigmoid_prime <= 5'b10001; end
				10'b0011010110: begin sigmoid <= 7'b1101100; sigmoid_prime <= 5'b10001; end
				10'b0011010111: begin sigmoid <= 7'b1101100; sigmoid_prime <= 5'b10001; end
				10'b0011011000: begin sigmoid <= 7'b1101100; sigmoid_prime <= 5'b10001; end
				10'b0011011001: begin sigmoid <= 7'b1101100; sigmoid_prime <= 5'b10001; end
				10'b0011011010: begin sigmoid <= 7'b1101100; sigmoid_prime <= 5'b10001; end
				10'b0011011011: begin sigmoid <= 7'b1101100; sigmoid_prime <= 5'b10001; end
				10'b0011011100: begin sigmoid <= 7'b1101101; sigmoid_prime <= 5'b10001; end
				10'b0011011101: begin sigmoid <= 7'b1101101; sigmoid_prime <= 5'b10000; end
				10'b0011011110: begin sigmoid <= 7'b1101101; sigmoid_prime <= 5'b10000; end
				10'b0011011111: begin sigmoid <= 7'b1101101; sigmoid_prime <= 5'b10000; end
				10'b0011100000: begin sigmoid <= 7'b1101101; sigmoid_prime <= 5'b10000; end
				10'b0011100001: begin sigmoid <= 7'b1101101; sigmoid_prime <= 5'b10000; end
				10'b0011100010: begin sigmoid <= 7'b1101101; sigmoid_prime <= 5'b10000; end
				10'b0011100011: begin sigmoid <= 7'b1101101; sigmoid_prime <= 5'b10000; end
				10'b0011100100: begin sigmoid <= 7'b1101110; sigmoid_prime <= 5'b10000; end
				10'b0011100101: begin sigmoid <= 7'b1101110; sigmoid_prime <= 5'b10000; end
				10'b0011100110: begin sigmoid <= 7'b1101110; sigmoid_prime <= 5'b10000; end
				10'b0011100111: begin sigmoid <= 7'b1101110; sigmoid_prime <= 5'b10000; end
				10'b0011101000: begin sigmoid <= 7'b1101110; sigmoid_prime <= 5'b01111; end
				10'b0011101001: begin sigmoid <= 7'b1101110; sigmoid_prime <= 5'b01111; end
				10'b0011101010: begin sigmoid <= 7'b1101110; sigmoid_prime <= 5'b01111; end
				10'b0011101011: begin sigmoid <= 7'b1101110; sigmoid_prime <= 5'b01111; end
				10'b0011101100: begin sigmoid <= 7'b1101111; sigmoid_prime <= 5'b01111; end
				10'b0011101101: begin sigmoid <= 7'b1101111; sigmoid_prime <= 5'b01111; end
				10'b0011101110: begin sigmoid <= 7'b1101111; sigmoid_prime <= 5'b01111; end
				10'b0011101111: begin sigmoid <= 7'b1101111; sigmoid_prime <= 5'b01111; end
				10'b0011110000: begin sigmoid <= 7'b1101111; sigmoid_prime <= 5'b01111; end
				10'b0011110001: begin sigmoid <= 7'b1101111; sigmoid_prime <= 5'b01111; end
				10'b0011110010: begin sigmoid <= 7'b1101111; sigmoid_prime <= 5'b01111; end
				10'b0011110011: begin sigmoid <= 7'b1101111; sigmoid_prime <= 5'b01111; end
				10'b0011110100: begin sigmoid <= 7'b1101111; sigmoid_prime <= 5'b01110; end
				10'b0011110101: begin sigmoid <= 7'b1110000; sigmoid_prime <= 5'b01110; end
				10'b0011110110: begin sigmoid <= 7'b1110000; sigmoid_prime <= 5'b01110; end
				10'b0011110111: begin sigmoid <= 7'b1110000; sigmoid_prime <= 5'b01110; end
				10'b0011111000: begin sigmoid <= 7'b1110000; sigmoid_prime <= 5'b01110; end
				10'b0011111001: begin sigmoid <= 7'b1110000; sigmoid_prime <= 5'b01110; end
				10'b0011111010: begin sigmoid <= 7'b1110000; sigmoid_prime <= 5'b01110; end
				10'b0011111011: begin sigmoid <= 7'b1110000; sigmoid_prime <= 5'b01110; end
				10'b0011111100: begin sigmoid <= 7'b1110000; sigmoid_prime <= 5'b01110; end
				10'b0011111101: begin sigmoid <= 7'b1110000; sigmoid_prime <= 5'b01110; end
				10'b0011111110: begin sigmoid <= 7'b1110001; sigmoid_prime <= 5'b01110; end
				10'b0011111111: begin sigmoid <= 7'b1110001; sigmoid_prime <= 5'b01110; end
				10'b0100000000: begin sigmoid <= 7'b1110001; sigmoid_prime <= 5'b01101; end
				10'b0100000001: begin sigmoid <= 7'b1110001; sigmoid_prime <= 5'b01101; end
				10'b0100000010: begin sigmoid <= 7'b1110001; sigmoid_prime <= 5'b01101; end
				10'b0100000011: begin sigmoid <= 7'b1110001; sigmoid_prime <= 5'b01101; end
				10'b0100000100: begin sigmoid <= 7'b1110001; sigmoid_prime <= 5'b01101; end
				10'b0100000101: begin sigmoid <= 7'b1110001; sigmoid_prime <= 5'b01101; end
				10'b0100000110: begin sigmoid <= 7'b1110001; sigmoid_prime <= 5'b01101; end
				10'b0100000111: begin sigmoid <= 7'b1110001; sigmoid_prime <= 5'b01101; end
				10'b0100001000: begin sigmoid <= 7'b1110010; sigmoid_prime <= 5'b01101; end
				10'b0100001001: begin sigmoid <= 7'b1110010; sigmoid_prime <= 5'b01101; end
				10'b0100001010: begin sigmoid <= 7'b1110010; sigmoid_prime <= 5'b01101; end
				10'b0100001011: begin sigmoid <= 7'b1110010; sigmoid_prime <= 5'b01101; end
				10'b0100001100: begin sigmoid <= 7'b1110010; sigmoid_prime <= 5'b01101; end
				10'b0100001101: begin sigmoid <= 7'b1110010; sigmoid_prime <= 5'b01100; end
				10'b0100001110: begin sigmoid <= 7'b1110010; sigmoid_prime <= 5'b01100; end
				10'b0100001111: begin sigmoid <= 7'b1110010; sigmoid_prime <= 5'b01100; end
				10'b0100010000: begin sigmoid <= 7'b1110010; sigmoid_prime <= 5'b01100; end
				10'b0100010001: begin sigmoid <= 7'b1110010; sigmoid_prime <= 5'b01100; end
				10'b0100010010: begin sigmoid <= 7'b1110011; sigmoid_prime <= 5'b01100; end
				10'b0100010011: begin sigmoid <= 7'b1110011; sigmoid_prime <= 5'b01100; end
				10'b0100010100: begin sigmoid <= 7'b1110011; sigmoid_prime <= 5'b01100; end
				10'b0100010101: begin sigmoid <= 7'b1110011; sigmoid_prime <= 5'b01100; end
				10'b0100010110: begin sigmoid <= 7'b1110011; sigmoid_prime <= 5'b01100; end
				10'b0100010111: begin sigmoid <= 7'b1110011; sigmoid_prime <= 5'b01100; end
				10'b0100011000: begin sigmoid <= 7'b1110011; sigmoid_prime <= 5'b01100; end
				10'b0100011001: begin sigmoid <= 7'b1110011; sigmoid_prime <= 5'b01100; end
				10'b0100011010: begin sigmoid <= 7'b1110011; sigmoid_prime <= 5'b01011; end
				10'b0100011011: begin sigmoid <= 7'b1110011; sigmoid_prime <= 5'b01011; end
				10'b0100011100: begin sigmoid <= 7'b1110011; sigmoid_prime <= 5'b01011; end
				10'b0100011101: begin sigmoid <= 7'b1110100; sigmoid_prime <= 5'b01011; end
				10'b0100011110: begin sigmoid <= 7'b1110100; sigmoid_prime <= 5'b01011; end
				10'b0100011111: begin sigmoid <= 7'b1110100; sigmoid_prime <= 5'b01011; end
				10'b0100100000: begin sigmoid <= 7'b1110100; sigmoid_prime <= 5'b01011; end
				10'b0100100001: begin sigmoid <= 7'b1110100; sigmoid_prime <= 5'b01011; end
				10'b0100100010: begin sigmoid <= 7'b1110100; sigmoid_prime <= 5'b01011; end
				10'b0100100011: begin sigmoid <= 7'b1110100; sigmoid_prime <= 5'b01011; end
				10'b0100100100: begin sigmoid <= 7'b1110100; sigmoid_prime <= 5'b01011; end
				10'b0100100101: begin sigmoid <= 7'b1110100; sigmoid_prime <= 5'b01011; end
				10'b0100100110: begin sigmoid <= 7'b1110100; sigmoid_prime <= 5'b01011; end
				10'b0100100111: begin sigmoid <= 7'b1110100; sigmoid_prime <= 5'b01011; end
				10'b0100101000: begin sigmoid <= 7'b1110100; sigmoid_prime <= 5'b01010; end
				10'b0100101001: begin sigmoid <= 7'b1110101; sigmoid_prime <= 5'b01010; end
				10'b0100101010: begin sigmoid <= 7'b1110101; sigmoid_prime <= 5'b01010; end
				10'b0100101011: begin sigmoid <= 7'b1110101; sigmoid_prime <= 5'b01010; end
				10'b0100101100: begin sigmoid <= 7'b1110101; sigmoid_prime <= 5'b01010; end
				10'b0100101101: begin sigmoid <= 7'b1110101; sigmoid_prime <= 5'b01010; end
				10'b0100101110: begin sigmoid <= 7'b1110101; sigmoid_prime <= 5'b01010; end
				10'b0100101111: begin sigmoid <= 7'b1110101; sigmoid_prime <= 5'b01010; end
				10'b0100110000: begin sigmoid <= 7'b1110101; sigmoid_prime <= 5'b01010; end
				10'b0100110001: begin sigmoid <= 7'b1110101; sigmoid_prime <= 5'b01010; end
				10'b0100110010: begin sigmoid <= 7'b1110101; sigmoid_prime <= 5'b01010; end
				10'b0100110011: begin sigmoid <= 7'b1110101; sigmoid_prime <= 5'b01010; end
				10'b0100110100: begin sigmoid <= 7'b1110101; sigmoid_prime <= 5'b01010; end
				10'b0100110101: begin sigmoid <= 7'b1110101; sigmoid_prime <= 5'b01010; end
				10'b0100110110: begin sigmoid <= 7'b1110110; sigmoid_prime <= 5'b01010; end
				10'b0100110111: begin sigmoid <= 7'b1110110; sigmoid_prime <= 5'b01010; end
				10'b0100111000: begin sigmoid <= 7'b1110110; sigmoid_prime <= 5'b01001; end
				10'b0100111001: begin sigmoid <= 7'b1110110; sigmoid_prime <= 5'b01001; end
				10'b0100111010: begin sigmoid <= 7'b1110110; sigmoid_prime <= 5'b01001; end
				10'b0100111011: begin sigmoid <= 7'b1110110; sigmoid_prime <= 5'b01001; end
				10'b0100111100: begin sigmoid <= 7'b1110110; sigmoid_prime <= 5'b01001; end
				10'b0100111101: begin sigmoid <= 7'b1110110; sigmoid_prime <= 5'b01001; end
				10'b0100111110: begin sigmoid <= 7'b1110110; sigmoid_prime <= 5'b01001; end
				10'b0100111111: begin sigmoid <= 7'b1110110; sigmoid_prime <= 5'b01001; end
				10'b0101000000: begin sigmoid <= 7'b1110110; sigmoid_prime <= 5'b01001; end
				10'b0101000001: begin sigmoid <= 7'b1110110; sigmoid_prime <= 5'b01001; end
				10'b0101000010: begin sigmoid <= 7'b1110110; sigmoid_prime <= 5'b01001; end
				10'b0101000011: begin sigmoid <= 7'b1110110; sigmoid_prime <= 5'b01001; end
				10'b0101000100: begin sigmoid <= 7'b1110111; sigmoid_prime <= 5'b01001; end
				10'b0101000101: begin sigmoid <= 7'b1110111; sigmoid_prime <= 5'b01001; end
				10'b0101000110: begin sigmoid <= 7'b1110111; sigmoid_prime <= 5'b01001; end
				10'b0101000111: begin sigmoid <= 7'b1110111; sigmoid_prime <= 5'b01001; end
				10'b0101001000: begin sigmoid <= 7'b1110111; sigmoid_prime <= 5'b01001; end
				10'b0101001001: begin sigmoid <= 7'b1110111; sigmoid_prime <= 5'b01000; end
				10'b0101001010: begin sigmoid <= 7'b1110111; sigmoid_prime <= 5'b01000; end
				10'b0101001011: begin sigmoid <= 7'b1110111; sigmoid_prime <= 5'b01000; end
				10'b0101001100: begin sigmoid <= 7'b1110111; sigmoid_prime <= 5'b01000; end
				10'b0101001101: begin sigmoid <= 7'b1110111; sigmoid_prime <= 5'b01000; end
				10'b0101001110: begin sigmoid <= 7'b1110111; sigmoid_prime <= 5'b01000; end
				10'b0101001111: begin sigmoid <= 7'b1110111; sigmoid_prime <= 5'b01000; end
				10'b0101010000: begin sigmoid <= 7'b1110111; sigmoid_prime <= 5'b01000; end
				10'b0101010001: begin sigmoid <= 7'b1110111; sigmoid_prime <= 5'b01000; end
				10'b0101010010: begin sigmoid <= 7'b1110111; sigmoid_prime <= 5'b01000; end
				10'b0101010011: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b01000; end
				10'b0101010100: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b01000; end
				10'b0101010101: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b01000; end
				10'b0101010110: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b01000; end
				10'b0101010111: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b01000; end
				10'b0101011000: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b01000; end
				10'b0101011001: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b01000; end
				10'b0101011010: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b01000; end
				10'b0101011011: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b00111; end
				10'b0101011100: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b00111; end
				10'b0101011101: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b00111; end
				10'b0101011110: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b00111; end
				10'b0101011111: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b00111; end
				10'b0101100000: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b00111; end
				10'b0101100001: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b00111; end
				10'b0101100010: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b00111; end
				10'b0101100011: begin sigmoid <= 7'b1111000; sigmoid_prime <= 5'b00111; end
				10'b0101100100: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00111; end
				10'b0101100101: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00111; end
				10'b0101100110: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00111; end
				10'b0101100111: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00111; end
				10'b0101101000: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00111; end
				10'b0101101001: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00111; end
				10'b0101101010: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00111; end
				10'b0101101011: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00111; end
				10'b0101101100: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00111; end
				10'b0101101101: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00111; end
				10'b0101101110: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00111; end
				10'b0101101111: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00111; end
				10'b0101110000: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00110; end
				10'b0101110001: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00110; end
				10'b0101110010: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00110; end
				10'b0101110011: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00110; end
				10'b0101110100: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00110; end
				10'b0101110101: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00110; end
				10'b0101110110: begin sigmoid <= 7'b1111001; sigmoid_prime <= 5'b00110; end
				10'b0101110111: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0101111000: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0101111001: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0101111010: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0101111011: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0101111100: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0101111101: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0101111110: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0101111111: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0110000000: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0110000001: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0110000010: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0110000011: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0110000100: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0110000101: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0110000110: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0110000111: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00110; end
				10'b0110001000: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00101; end
				10'b0110001001: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00101; end
				10'b0110001010: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00101; end
				10'b0110001011: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00101; end
				10'b0110001100: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00101; end
				10'b0110001101: begin sigmoid <= 7'b1111010; sigmoid_prime <= 5'b00101; end
				10'b0110001110: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110001111: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110010000: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110010001: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110010010: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110010011: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110010100: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110010101: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110010110: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110010111: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110011000: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110011001: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110011010: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110011011: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110011100: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110011101: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110011110: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110011111: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110100000: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110100001: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110100010: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110100011: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00101; end
				10'b0110100100: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00100; end
				10'b0110100101: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00100; end
				10'b0110100110: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00100; end
				10'b0110100111: begin sigmoid <= 7'b1111011; sigmoid_prime <= 5'b00100; end
				10'b0110101000: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110101001: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110101010: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110101011: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110101100: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110101101: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110101110: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110101111: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110110000: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110110001: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110110010: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110110011: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110110100: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110110101: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110110110: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110110111: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110111000: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110111001: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110111010: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110111011: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110111100: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110111101: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110111110: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0110111111: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0111000000: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0111000001: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0111000010: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0111000011: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0111000100: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0111000101: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00100; end
				10'b0111000110: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00011; end
				10'b0111000111: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00011; end
				10'b0111001000: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00011; end
				10'b0111001001: begin sigmoid <= 7'b1111100; sigmoid_prime <= 5'b00011; end
				10'b0111001010: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111001011: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111001100: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111001101: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111001110: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111001111: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111010000: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111010001: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111010010: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111010011: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111010100: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111010101: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111010110: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111010111: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111011000: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111011001: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111011010: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111011011: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111011100: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111011101: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111011110: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111011111: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111100000: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111100001: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111100010: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111100011: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111100100: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111100101: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111100110: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111100111: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111101000: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111101001: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111101010: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111101011: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111101100: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111101101: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111101110: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111101111: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111110000: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111110001: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111110010: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00011; end
				10'b0111110011: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00010; end
				10'b0111110100: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00010; end
				10'b0111110101: begin sigmoid <= 7'b1111101; sigmoid_prime <= 5'b00010; end
				10'b0111110110: begin sigmoid <= 7'b1111110; sigmoid_prime <= 5'b00010; end
				10'b0111110111: begin sigmoid <= 7'b1111110; sigmoid_prime <= 5'b00010; end
				10'b0111111000: begin sigmoid <= 7'b1111110; sigmoid_prime <= 5'b00010; end
				10'b0111111001: begin sigmoid <= 7'b1111110; sigmoid_prime <= 5'b00010; end
				10'b0111111010: begin sigmoid <= 7'b1111110; sigmoid_prime <= 5'b00010; end
				10'b0111111011: begin sigmoid <= 7'b1111110; sigmoid_prime <= 5'b00010; end
				10'b0111111100: begin sigmoid <= 7'b1111110; sigmoid_prime <= 5'b00010; end
				10'b0111111101: begin sigmoid <= 7'b1111110; sigmoid_prime <= 5'b00010; end
				10'b0111111110: begin sigmoid <= 7'b1111110; sigmoid_prime <= 5'b00010; end
				10'b0111111111: begin sigmoid <= 7'b1111110; sigmoid_prime <= 5'b00010; end
		
	endcase
	end
endmodule
